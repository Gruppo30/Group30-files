LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.ALL;

entity InstructionMemory is
	generic ( 	k : positive := 8);
	port(	clk,rst     : in std_logic;
			addr 	   : in  std_logic_vector(31 downto 0);
			data_out   : out std_logic_vector(31 downto 0)
		);
end InstructionMemory;

architecture beh of InstructionMemory is

	type mem is array(0 to (2**k)-1)  of std_logic_vector (31 downto 0);
	signal memArray : mem := (others => "00000000000000000000000000000000");
				
begin 

	memArray(0 to 31) <= (		"00000000011100000000100000010011",
								"00001111110000010000001000010111",
								"11111111110000100000001000010011",
								"00001111110000010000001010010111",
								"00000001000000101000001010010011",
								"01000000000000000000011010110111",
								"11111111111101101000011010010011",
								"00000010000010000000001001100011",
								"00000000000000100010010000000011",
								"00000000000001000000010100100111",
								"00000000010000100000001000010011",
								"11111111111110000000100000010011",
								"00000000110101010010010110110011",
								"11111110000001011000010011100011",
								"00000000000001010000011010110011",
								"11111110000111111111000011101111",
								"00000000110100101010000000100011",
								"00000000000000000000000000010011",
								"00000000000000000000000000000000",
								"00000000000000000000000000000000",
								"00000000000000000000000000000000",
								"00000000000000000000000000000000",
								"00000000000000000000000000000000",
								"00000000000000000000000000000000",
								"00000000000000000000000000000000",
								"00000000000000000000000000000000",
								"00000000000000000000000000000000",
								"00000000000000000000000000000000",
								"00000000000000000000000000000000",
								"00000000000000000000000000000000",
								"00000000000000000000000000000000",
								"00000000000000000000000000000000");

	process(addr, rst) is
	begin
		if(rst = '0') then
--			data_out <= (others => '0');
			data_out <= memArray(0);
		else
			data_out <= memArray((to_integer(unsigned(addr(7 downto 0))))/4);
		end if;
	end process;

end beh;

