library ieee;
use ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

-- This file has been automatically generated though the C code which can be found 
-- in the appendix of the lab reports. We are not going to comment it since it is 
-- just a connection and a series of instances of HA and FA components 
-- useful to implement the dadda tree

entity dadda_tree is
	port (y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17 : in std_logic_vector (63 downto 0);
			product : OUT std_logic_vector(63 downto 0)
		  );
end dadda_tree;

architecture beh of dadda_tree is

component FA is
port ( a_fa, b_fa, cin_fa : IN std_logic;
	s_fa, c_fa : OUT std_logic);
end component fa;

component HA is
port ( a_ha, b_ha : IN std_logic;
	s_ha, c_ha : OUT std_logic);
end component ha;
	
	signal p0_y0,p0_y1,p0_y2,p0_y3,p0_y4,p0_y5,p0_y6,p0_y7,p0_y8,p0_y9,p0_y10,p0_y11,p0_y12,p0_y13,p0_y14,p0_y15,p0_y16 : std_logic_vector (63 downto 0);
	signal p1_y0,p1_y1,p1_y2,p1_y3,p1_y4,p1_y5,p1_y6,p1_y7,p1_y8,p1_y9,p1_y10,p1_y11,p1_y12 : std_logic_vector (63 downto 0);
	signal p2_y0,p2_y1,p2_y2,p2_y3,p2_y4,p2_y5,p2_y6,p2_y7,p2_y8 : std_logic_vector (63 downto 0);
	signal p3_y0,p3_y1,p3_y2,p3_y3,p3_y4,p3_y5 : std_logic_vector (63 downto 0);
	signal p4_y0,p4_y1,p4_y2,p4_y3 : std_logic_vector (63 downto 0);
	signal p5_y0,p5_y1,p5_y2 : std_logic_vector (63 downto 0);
	signal p6_y0,p6_y1 : std_logic_vector (63 downto 0);
	signal overflow_bit: std_logic;
	
begin

	p0_y0<=y16(63)&y15(62 downto 61)&y14(60 downto 59)&y13(58 downto 57)&y12(56 downto 55)&y11(54 downto 53)&y10(52 downto 51)&y9(50 downto 49)&y8(48 downto 47)&y7(46 downto 45)&y6(44 downto 43)&y5(42 downto 41)&y4(40 downto 39)&y3(38 downto 37)&y2(36)&y1(35 downto 0);
	p0_y1<=y17(63)&y16(62 downto 61)&y15(60 downto 59)&y14(58 downto 57)&y13(56 downto 55)&y12(54 downto 53)&y11(52 downto 51)&y10(50 downto 49)&y9(48 downto 47)&y8(46 downto 45)&y7(44 downto 43)&y6(42 downto 41)&y5(40 downto 39)&y4(38 downto 37)&y3(36)&y2(35 downto 0);
	p0_y2<='Z'&y17(62 downto 61)&y16(60 downto 59)&y15(58 downto 57)&y14(56 downto 55)&y13(54 downto 53)&y12(52 downto 51)&y11(50 downto 49)&y10(48 downto 47)&y9(46 downto 45)&y8(44 downto 43)&y7(42 downto 41)&y6(40 downto 39)&y5(38 downto 37)&y4(36)&y3(35 downto 0);
	p0_y3<="ZZZ"&y17(60 downto 59)&y16(58 downto 57)&y15(56 downto 55)&y14(54 downto 53)&y13(52 downto 51)&y12(50 downto 49)&y11(48 downto 47)&y10(46 downto 45)&y9(44 downto 43)&y8(42 downto 41)&y7(40 downto 39)&y6(38 downto 37)&y5(36)&y4(35 downto 0);
	p0_y4<="ZZZZZ"&y17(58 downto 57)&y16(56 downto 55)&y15(54 downto 53)&y14(52 downto 51)&y13(50 downto 49)&y12(48 downto 47)&y11(46 downto 45)&y10(44 downto 43)&y9(42 downto 41)&y8(40 downto 39)&y7(38 downto 37)&y6(36)&y5(35 downto 0);
	p0_y5<="ZZZZZZZ"&y17(56 downto 55)&y16(54 downto 53)&y15(52 downto 51)&y14(50 downto 49)&y13(48 downto 47)&y12(46 downto 45)&y11(44 downto 43)&y10(42 downto 41)&y9(40 downto 39)&y8(38 downto 37)&y7(36)&y6(35 downto 0);
	p0_y6<="ZZZZZZZZZ"&y17(54 downto 53)&y16(52 downto 51)&y15(50 downto 49)&y14(48 downto 47)&y13(46 downto 45)&y12(44 downto 43)&y11(42 downto 41)&y10(40 downto 39)&y9(38 downto 37)&y8(36)&y7(35 downto 0);
	p0_y7<="ZZZZZZZZZZZ"&y17(52 downto 51)&y16(50 downto 49)&y15(48 downto 47)&y14(46 downto 45)&y13(44 downto 43)&y12(42 downto 41)&y11(40 downto 39)&y10(38 downto 37)&y9(36)&y8(35 downto 0);
	p0_y8<="ZZZZZZZZZZZZZ"&y17(50 downto 49)&y16(48 downto 47)&y15(46 downto 45)&y14(44 downto 43)&y13(42 downto 41)&y12(40 downto 39)&y11(38 downto 37)&y10(36)&y9(35 downto 0);
	p0_y9<="ZZZZZZZZZZZZZZZ"&y17(48 downto 47)&y16(46 downto 45)&y15(44 downto 43)&y14(42 downto 41)&y13(40 downto 39)&y12(38 downto 37)&y11(36)&y10(35 downto 0);
	p0_y10<="ZZZZZZZZZZZZZZZZZ"&y17(46 downto 45)&y16(44 downto 43)&y15(42 downto 41)&y14(40 downto 39)&y13(38 downto 37)&y12(36)&y11(35 downto 0);
	p0_y11<="ZZZZZZZZZZZZZZZZZZZ"&y17(44 downto 43)&y16(42 downto 41)&y15(40 downto 39)&y14(38 downto 37)&y13(36)&y12(35 downto 0);
	p0_y12<="ZZZZZZZZZZZZZZZZZZZZZ"&y17(42 downto 41)&y16(40 downto 39)&y15(38 downto 37)&y14(36)&y13(35 downto 0);
	p0_y13<="ZZZZZZZZZZZZZZZZZZZZZZZ"&y17(40 downto 39)&y16(38 downto 37)&y15(36)&y14(35 downto 0);
	p0_y14<="ZZZZZZZZZZZZZZZZZZZZZZZZZ"&y17(38 downto 37)&y16(36)&y15(35 downto 0);
	p0_y15<="ZZZZZZZZZZZZZZZZZZZZZZZZZZZ"&y17(36)&y16(35 downto 0);
	p0_y16<="ZZZZZZZZZZZZZZZZZZZZZZZZZZZZ"&y16(35 downto 0);
	
	p1_y0(0)<=p0_y0(0);
	p1_y1(0)<=p0_y1(0);
	p1_y0(1)<=p0_y0(1);
	p1_y1(1)<=p0_y1(1);
	p1_y0(2)<=p0_y0(2);
	p1_y1(2)<=p0_y1(2);
	p1_y2(2)<=p0_y2(2);
	p1_y0(3)<=p0_y0(3);
	p1_y1(3)<=p0_y1(3);
	p1_y2(3)<=p0_y2(3);
	p1_y0(4)<=p0_y0(4);
	p1_y1(4)<=p0_y1(4);
	p1_y2(4)<=p0_y2(4);
	p1_y3(4)<=p0_y3(4);
	p1_y0(5)<=p0_y0(5);
	p1_y1(5)<=p0_y1(5);
	p1_y2(5)<=p0_y2(5);
	p1_y3(5)<=p0_y3(5);
	p1_y0(6)<=p0_y0(6);
	p1_y1(6)<=p0_y1(6);
	p1_y2(6)<=p0_y2(6);
	p1_y3(6)<=p0_y3(6);
	p1_y4(6)<=p0_y4(6);
	p1_y0(7)<=p0_y0(7);
	p1_y1(7)<=p0_y1(7);
	p1_y2(7)<=p0_y2(7);
	p1_y3(7)<=p0_y3(7);
	p1_y4(7)<=p0_y4(7);
	p1_y0(8)<=p0_y0(8);
	p1_y1(8)<=p0_y1(8);
	p1_y2(8)<=p0_y2(8);
	p1_y3(8)<=p0_y3(8);
	p1_y4(8)<=p0_y4(8);
	p1_y5(8)<=p0_y5(8);
	p1_y0(9)<=p0_y0(9);
	p1_y1(9)<=p0_y1(9);
	p1_y2(9)<=p0_y2(9);
	p1_y3(9)<=p0_y3(9);
	p1_y4(9)<=p0_y4(9);
	p1_y5(9)<=p0_y5(9);
	p1_y0(10)<=p0_y0(10);
	p1_y1(10)<=p0_y1(10);
	p1_y2(10)<=p0_y2(10);
	p1_y3(10)<=p0_y3(10);
	p1_y4(10)<=p0_y4(10);
	p1_y5(10)<=p0_y5(10);
	p1_y6(10)<=p0_y6(10);
	p1_y0(11)<=p0_y0(11);
	p1_y1(11)<=p0_y1(11);
	p1_y2(11)<=p0_y2(11);
	p1_y3(11)<=p0_y3(11);
	p1_y4(11)<=p0_y4(11);
	p1_y5(11)<=p0_y5(11);
	p1_y6(11)<=p0_y6(11);
	p1_y0(12)<=p0_y0(12);
	p1_y1(12)<=p0_y1(12);
	p1_y2(12)<=p0_y2(12);
	p1_y3(12)<=p0_y3(12);
	p1_y4(12)<=p0_y4(12);
	p1_y5(12)<=p0_y5(12);
	p1_y6(12)<=p0_y6(12);
	p1_y7(12)<=p0_y7(12);
	p1_y0(13)<=p0_y0(13);
	p1_y1(13)<=p0_y1(13);
	p1_y2(13)<=p0_y2(13);
	p1_y3(13)<=p0_y3(13);
	p1_y4(13)<=p0_y4(13);
	p1_y5(13)<=p0_y5(13);
	p1_y6(13)<=p0_y6(13);
	p1_y7(13)<=p0_y7(13);
	p1_y0(14)<=p0_y0(14);
	p1_y1(14)<=p0_y1(14);
	p1_y2(14)<=p0_y2(14);
	p1_y3(14)<=p0_y3(14);
	p1_y4(14)<=p0_y4(14);
	p1_y5(14)<=p0_y5(14);
	p1_y6(14)<=p0_y6(14);
	p1_y7(14)<=p0_y7(14);
	p1_y8(14)<=p0_y8(14);
	p1_y0(15)<=p0_y0(15);
	p1_y1(15)<=p0_y1(15);
	p1_y2(15)<=p0_y2(15);
	p1_y3(15)<=p0_y3(15);
	p1_y4(15)<=p0_y4(15);
	p1_y5(15)<=p0_y5(15);
	p1_y6(15)<=p0_y6(15);
	p1_y7(15)<=p0_y7(15);
	p1_y8(15)<=p0_y8(15);
	p1_y0(16)<=p0_y0(16);
	p1_y1(16)<=p0_y1(16);
	p1_y2(16)<=p0_y2(16);
	p1_y3(16)<=p0_y3(16);
	p1_y4(16)<=p0_y4(16);
	p1_y5(16)<=p0_y5(16);
	p1_y6(16)<=p0_y6(16);
	p1_y7(16)<=p0_y7(16);
	p1_y8(16)<=p0_y8(16);
	p1_y9(16)<=p0_y9(16);
	p1_y0(17)<=p0_y0(17);
	p1_y1(17)<=p0_y1(17);
	p1_y2(17)<=p0_y2(17);
	p1_y3(17)<=p0_y3(17);
	p1_y4(17)<=p0_y4(17);
	p1_y5(17)<=p0_y5(17);
	p1_y6(17)<=p0_y6(17);
	p1_y7(17)<=p0_y7(17);
	p1_y8(17)<=p0_y8(17);
	p1_y9(17)<=p0_y9(17);
	p1_y0(18)<=p0_y0(18);
	p1_y1(18)<=p0_y1(18);
	p1_y2(18)<=p0_y2(18);
	p1_y3(18)<=p0_y3(18);
	p1_y4(18)<=p0_y4(18);
	p1_y5(18)<=p0_y5(18);
	p1_y6(18)<=p0_y6(18);
	p1_y7(18)<=p0_y7(18);
	p1_y8(18)<=p0_y8(18);
	p1_y9(18)<=p0_y9(18);
	p1_y10(18)<=p0_y10(18);
	p1_y0(19)<=p0_y0(19);
	p1_y1(19)<=p0_y1(19);
	p1_y2(19)<=p0_y2(19);
	p1_y3(19)<=p0_y3(19);
	p1_y4(19)<=p0_y4(19);
	p1_y5(19)<=p0_y5(19);
	p1_y6(19)<=p0_y6(19);
	p1_y7(19)<=p0_y7(19);
	p1_y8(19)<=p0_y8(19);
	p1_y9(19)<=p0_y9(19);
	p1_y10(19)<=p0_y10(19);
	p1_y0(20)<=p0_y0(20);
	p1_y1(20)<=p0_y1(20);
	p1_y2(20)<=p0_y2(20);
	p1_y3(20)<=p0_y3(20);
	p1_y4(20)<=p0_y4(20);
	p1_y5(20)<=p0_y5(20);
	p1_y6(20)<=p0_y6(20);
	p1_y7(20)<=p0_y7(20);
	p1_y8(20)<=p0_y8(20);
	p1_y9(20)<=p0_y9(20);
	p1_y10(20)<=p0_y10(20);
	p1_y11(20)<=p0_y11(20);
	p1_y0(21)<=p0_y0(21);
	p1_y1(21)<=p0_y1(21);
	p1_y2(21)<=p0_y2(21);
	p1_y3(21)<=p0_y3(21);
	p1_y4(21)<=p0_y4(21);
	p1_y5(21)<=p0_y5(21);
	p1_y6(21)<=p0_y6(21);
	p1_y7(21)<=p0_y7(21);
	p1_y8(21)<=p0_y8(21);
	p1_y9(21)<=p0_y9(21);
	p1_y10(21)<=p0_y10(21);
	p1_y11(21)<=p0_y11(21);
	p1_y0(22)<=p0_y0(22);
	p1_y1(22)<=p0_y1(22);
	p1_y2(22)<=p0_y2(22);
	p1_y3(22)<=p0_y3(22);
	p1_y4(22)<=p0_y4(22);
	p1_y5(22)<=p0_y5(22);
	p1_y6(22)<=p0_y6(22);
	p1_y7(22)<=p0_y7(22);
	p1_y8(22)<=p0_y8(22);
	p1_y9(22)<=p0_y9(22);
	p1_y10(22)<=p0_y10(22);
	p1_y11(22)<=p0_y11(22);
	p1_y12(22)<=p0_y12(22);
	p1_y0(23)<=p0_y0(23);
	p1_y1(23)<=p0_y1(23);
	p1_y2(23)<=p0_y2(23);
	p1_y3(23)<=p0_y3(23);
	p1_y4(23)<=p0_y4(23);
	p1_y5(23)<=p0_y5(23);
	p1_y6(23)<=p0_y6(23);
	p1_y7(23)<=p0_y7(23);
	p1_y8(23)<=p0_y8(23);
	p1_y9(23)<=p0_y9(23);
	p1_y10(23)<=p0_y10(23);
	p1_y11(23)<=p0_y11(23);
	p1_y12(23)<=p0_y12(23);
	HA0: HA PORT MAP (p0_y0(24),p0_y1(24),p1_y0(24),p1_y0(25));
	p1_y1(24)<=p0_y2(24);
	p1_y2(24)<=p0_y3(24);
	p1_y3(24)<=p0_y4(24);
	p1_y4(24)<=p0_y5(24);
	p1_y5(24)<=p0_y6(24);
	p1_y6(24)<=p0_y7(24);
	p1_y7(24)<=p0_y8(24);
	p1_y8(24)<=p0_y9(24);
	p1_y9(24)<=p0_y10(24);
	p1_y10(24)<=p0_y11(24);
	p1_y11(24)<=p0_y12(24);
	p1_y12(24)<=p0_y13(24);
	FA0: FA PORT MAP (p0_y0(25),p0_y1(25),p0_y2(25),p1_y1(25),p1_y0(26));
	p1_y2(25)<=p0_y3(25);
	p1_y3(25)<=p0_y4(25);
	p1_y4(25)<=p0_y5(25);
	p1_y5(25)<=p0_y6(25);
	p1_y6(25)<=p0_y7(25);
	p1_y7(25)<=p0_y8(25);
	p1_y8(25)<=p0_y9(25);
	p1_y9(25)<=p0_y10(25);
	p1_y10(25)<=p0_y11(25);
	p1_y11(25)<=p0_y12(25);
	p1_y12(25)<=p0_y13(25);
	FA1: FA PORT MAP (p0_y0(26),p0_y1(26),p0_y2(26),p1_y1(26),p1_y0(27));
	HA1: HA PORT MAP (p0_y3(26),p0_y4(26),p1_y2(26),p1_y1(27));
	p1_y3(26)<=p0_y5(26);
	p1_y4(26)<=p0_y6(26);
	p1_y5(26)<=p0_y7(26);
	p1_y6(26)<=p0_y8(26);
	p1_y7(26)<=p0_y9(26);
	p1_y8(26)<=p0_y10(26);
	p1_y9(26)<=p0_y11(26);
	p1_y10(26)<=p0_y12(26);
	p1_y11(26)<=p0_y13(26);
	p1_y12(26)<=p0_y14(26);
	FA2: FA PORT MAP (p0_y0(27),p0_y1(27),p0_y2(27),p1_y2(27),p1_y0(28));
	FA3: FA PORT MAP (p0_y3(27),p0_y4(27),p0_y5(27),p1_y3(27),p1_y1(28));
	p1_y4(27)<=p0_y6(27);
	p1_y5(27)<=p0_y7(27);
	p1_y6(27)<=p0_y8(27);
	p1_y7(27)<=p0_y9(27);
	p1_y8(27)<=p0_y10(27);
	p1_y9(27)<=p0_y11(27);
	p1_y10(27)<=p0_y12(27);
	p1_y11(27)<=p0_y13(27);
	p1_y12(27)<=p0_y14(27);
	FA4: FA PORT MAP (p0_y0(28),p0_y1(28),p0_y2(28),p1_y2(28),p1_y0(29));
	FA5: FA PORT MAP (p0_y3(28),p0_y4(28),p0_y5(28),p1_y3(28),p1_y1(29));
	HA2: HA PORT MAP (p0_y6(28),p0_y7(28),p1_y4(28),p1_y2(29));
	p1_y5(28)<=p0_y8(28);
	p1_y6(28)<=p0_y9(28);
	p1_y7(28)<=p0_y10(28);
	p1_y8(28)<=p0_y11(28);
	p1_y9(28)<=p0_y12(28);
	p1_y10(28)<=p0_y13(28);
	p1_y11(28)<=p0_y14(28);
	p1_y12(28)<=p0_y15(28);
	FA6: FA PORT MAP (p0_y0(29),p0_y1(29),p0_y2(29),p1_y3(29),p1_y0(30));
	FA7: FA PORT MAP (p0_y3(29),p0_y4(29),p0_y5(29),p1_y4(29),p1_y1(30));
	FA8: FA PORT MAP (p0_y6(29),p0_y7(29),p0_y8(29),p1_y5(29),p1_y2(30));
	p1_y6(29)<=p0_y9(29);
	p1_y7(29)<=p0_y10(29);
	p1_y8(29)<=p0_y11(29);
	p1_y9(29)<=p0_y12(29);
	p1_y10(29)<=p0_y13(29);
	p1_y11(29)<=p0_y14(29);
	p1_y12(29)<=p0_y15(29);
	FA9: FA PORT MAP (p0_y0(30),p0_y1(30),p0_y2(30),p1_y3(30),p1_y0(31));
	FA10: FA PORT MAP (p0_y3(30),p0_y4(30),p0_y5(30),p1_y4(30),p1_y1(31));
	FA11: FA PORT MAP (p0_y6(30),p0_y7(30),p0_y8(30),p1_y5(30),p1_y2(31));
	HA3: HA PORT MAP (p0_y9(30),p0_y10(30),p1_y6(30),p1_y3(31));
	p1_y7(30)<=p0_y11(30);
	p1_y8(30)<=p0_y12(30);
	p1_y9(30)<=p0_y13(30);
	p1_y10(30)<=p0_y14(30);
	p1_y11(30)<=p0_y15(30);
	p1_y12(30)<=p0_y16(30);
	FA12: FA PORT MAP (p0_y0(31),p0_y1(31),p0_y2(31),p1_y4(31),p1_y0(32));
	FA13: FA PORT MAP (p0_y3(31),p0_y4(31),p0_y5(31),p1_y5(31),p1_y1(32));
	FA14: FA PORT MAP (p0_y6(31),p0_y7(31),p0_y8(31),p1_y6(31),p1_y2(32));
	FA15: FA PORT MAP (p0_y9(31),p0_y10(31),p0_y11(31),p1_y7(31),p1_y3(32));
	p1_y8(31)<=p0_y12(31);
	p1_y9(31)<=p0_y13(31);
	p1_y10(31)<=p0_y14(31);
	p1_y11(31)<=p0_y15(31);
	p1_y12(31)<=p0_y16(31);
	FA16: FA PORT MAP (p0_y0(32),p0_y1(32),p0_y2(32),p1_y4(32),p1_y0(33));
	FA17: FA PORT MAP (p0_y3(32),p0_y4(32),p0_y5(32),p1_y5(32),p1_y1(33));
	FA18: FA PORT MAP (p0_y6(32),p0_y7(32),p0_y8(32),p1_y6(32),p1_y2(33));
	FA19: FA PORT MAP (p0_y9(32),p0_y10(32),p0_y11(32),p1_y7(32),p1_y3(33));
	p1_y8(32)<=p0_y12(32);
	p1_y9(32)<=p0_y13(32);
	p1_y10(32)<=p0_y14(32);
	p1_y11(32)<=p0_y15(32);
	p1_y12(32)<=p0_y16(32);
	FA20: FA PORT MAP (p0_y0(33),p0_y1(33),p0_y2(33),p1_y4(33),p1_y0(34));
	FA21: FA PORT MAP (p0_y3(33),p0_y4(33),p0_y5(33),p1_y5(33),p1_y1(34));
	FA22: FA PORT MAP (p0_y6(33),p0_y7(33),p0_y8(33),p1_y6(33),p1_y2(34));
	FA23: FA PORT MAP (p0_y9(33),p0_y10(33),p0_y11(33),p1_y7(33),p1_y3(34));
	p1_y8(33)<=p0_y12(33);
	p1_y9(33)<=p0_y13(33);
	p1_y10(33)<=p0_y14(33);
	p1_y11(33)<=p0_y15(33);
	p1_y12(33)<=p0_y16(33);
	FA24: FA PORT MAP (p0_y0(34),p0_y1(34),p0_y2(34),p1_y4(34),p1_y0(35));
	FA25: FA PORT MAP (p0_y3(34),p0_y4(34),p0_y5(34),p1_y5(34),p1_y1(35));
	FA26: FA PORT MAP (p0_y6(34),p0_y7(34),p0_y8(34),p1_y6(34),p1_y2(35));
	FA27: FA PORT MAP (p0_y9(34),p0_y10(34),p0_y11(34),p1_y7(34),p1_y3(35));
	p1_y8(34)<=p0_y12(34);
	p1_y9(34)<=p0_y13(34);
	p1_y10(34)<=p0_y14(34);
	p1_y11(34)<=p0_y15(34);
	p1_y12(34)<=p0_y16(34);
	FA28: FA PORT MAP (p0_y0(35),p0_y1(35),p0_y2(35),p1_y4(35),p1_y0(36));
	FA29: FA PORT MAP (p0_y3(35),p0_y4(35),p0_y5(35),p1_y5(35),p1_y1(36));
	FA30: FA PORT MAP (p0_y6(35),p0_y7(35),p0_y8(35),p1_y6(35),p1_y2(36));
	FA31: FA PORT MAP (p0_y9(35),p0_y10(35),p0_y11(35),p1_y7(35),p1_y3(36));
	p1_y8(35)<=p0_y12(35);
	p1_y9(35)<=p0_y13(35);
	p1_y10(35)<=p0_y14(35);
	p1_y11(35)<=p0_y15(35);
	p1_y12(35)<=p0_y16(35);
	FA32: FA PORT MAP (p0_y0(36),p0_y1(36),p0_y2(36),p1_y4(36),p1_y0(37));
	FA33: FA PORT MAP (p0_y3(36),p0_y4(36),p0_y5(36),p1_y5(36),p1_y1(37));
	FA34: FA PORT MAP (p0_y6(36),p0_y7(36),p0_y8(36),p1_y6(36),p1_y2(37));
	HA4: HA PORT MAP (p0_y9(36),p0_y10(36),p1_y7(36),p1_y3(37));
	p1_y8(36)<=p0_y11(36);
	p1_y9(36)<=p0_y12(36);
	p1_y10(36)<=p0_y13(36);
	p1_y11(36)<=p0_y14(36);
	p1_y12(36)<=p0_y15(36);
	FA35: FA PORT MAP (p0_y0(37),p0_y1(37),p0_y2(37),p1_y4(37),p1_y0(38));
	FA36: FA PORT MAP (p0_y3(37),p0_y4(37),p0_y5(37),p1_y5(37),p1_y1(38));
	FA37: FA PORT MAP (p0_y6(37),p0_y7(37),p0_y8(37),p1_y6(37),p1_y2(38));
	p1_y7(37)<=p0_y9(37);
	p1_y8(37)<=p0_y10(37);
	p1_y9(37)<=p0_y11(37);
	p1_y10(37)<=p0_y12(37);
	p1_y11(37)<=p0_y13(37);
	p1_y12(37)<=p0_y14(37);
	FA38: FA PORT MAP (p0_y0(38),p0_y1(38),p0_y2(38),p1_y3(38),p1_y0(39));
	FA39: FA PORT MAP (p0_y3(38),p0_y4(38),p0_y5(38),p1_y4(38),p1_y1(39));
	HA5: HA PORT MAP (p0_y6(38),p0_y7(38),p1_y5(38),p1_y2(39));
	p1_y6(38)<=p0_y8(38);
	p1_y7(38)<=p0_y9(38);
	p1_y8(38)<=p0_y10(38);
	p1_y9(38)<=p0_y11(38);
	p1_y10(38)<=p0_y12(38);
	p1_y11(38)<=p0_y13(38);
	p1_y12(38)<=p0_y14(38);
	FA40: FA PORT MAP (p0_y0(39),p0_y1(39),p0_y2(39),p1_y3(39),p1_y0(40));
	FA41: FA PORT MAP (p0_y3(39),p0_y4(39),p0_y5(39),p1_y4(39),p1_y1(40));
	p1_y5(39)<=p0_y6(39);
	p1_y6(39)<=p0_y7(39);
	p1_y7(39)<=p0_y8(39);
	p1_y8(39)<=p0_y9(39);
	p1_y9(39)<=p0_y10(39);
	p1_y10(39)<=p0_y11(39);
	p1_y11(39)<=p0_y12(39);
	p1_y12(39)<=p0_y13(39);
	FA42: FA PORT MAP (p0_y0(40),p0_y1(40),p0_y2(40),p1_y2(40),p1_y0(41));
	HA6: HA PORT MAP (p0_y3(40),p0_y4(40),p1_y3(40),p1_y1(41));
	p1_y4(40)<=p0_y5(40);
	p1_y5(40)<=p0_y6(40);
	p1_y6(40)<=p0_y7(40);
	p1_y7(40)<=p0_y8(40);
	p1_y8(40)<=p0_y9(40);
	p1_y9(40)<=p0_y10(40);
	p1_y10(40)<=p0_y11(40);
	p1_y11(40)<=p0_y12(40);
	p1_y12(40)<=p0_y13(40);
	FA43: FA PORT MAP (p0_y0(41),p0_y1(41),p0_y2(41),p1_y2(41),p1_y0(42));
	p1_y3(41)<=p0_y3(41);
	p1_y4(41)<=p0_y4(41);
	p1_y5(41)<=p0_y5(41);
	p1_y6(41)<=p0_y6(41);
	p1_y7(41)<=p0_y7(41);
	p1_y8(41)<=p0_y8(41);
	p1_y9(41)<=p0_y9(41);
	p1_y10(41)<=p0_y10(41);
	p1_y11(41)<=p0_y11(41);
	p1_y12(41)<=p0_y12(41);
	HA7: HA PORT MAP (p0_y0(42),p0_y1(42),p1_y1(42),p1_y0(43));
	p1_y2(42)<=p0_y2(42);
	p1_y3(42)<=p0_y3(42);
	p1_y4(42)<=p0_y4(42);
	p1_y5(42)<=p0_y5(42);
	p1_y6(42)<=p0_y6(42);
	p1_y7(42)<=p0_y7(42);
	p1_y8(42)<=p0_y8(42);
	p1_y9(42)<=p0_y9(42);
	p1_y10(42)<=p0_y10(42);
	p1_y11(42)<=p0_y11(42);
	p1_y12(42)<=p0_y12(42);
	p1_y1(43)<=p0_y0(43);
	p1_y2(43)<=p0_y1(43);
	p1_y3(43)<=p0_y2(43);
	p1_y4(43)<=p0_y3(43);
	p1_y5(43)<=p0_y4(43);
	p1_y6(43)<=p0_y5(43);
	p1_y7(43)<=p0_y6(43);
	p1_y8(43)<=p0_y7(43);
	p1_y9(43)<=p0_y8(43);
	p1_y10(43)<=p0_y9(43);
	p1_y11(43)<=p0_y10(43);
	p1_y12(43)<=p0_y11(43);
	p1_y0(44)<=p0_y0(44);
	p1_y1(44)<=p0_y1(44);
	p1_y2(44)<=p0_y2(44);
	p1_y3(44)<=p0_y3(44);
	p1_y4(44)<=p0_y4(44);
	p1_y5(44)<=p0_y5(44);
	p1_y6(44)<=p0_y6(44);
	p1_y7(44)<=p0_y7(44);
	p1_y8(44)<=p0_y8(44);
	p1_y9(44)<=p0_y9(44);
	p1_y10(44)<=p0_y10(44);
	p1_y11(44)<=p0_y11(44);
	p1_y0(45)<=p0_y0(45);
	p1_y1(45)<=p0_y1(45);
	p1_y2(45)<=p0_y2(45);
	p1_y3(45)<=p0_y3(45);
	p1_y4(45)<=p0_y4(45);
	p1_y5(45)<=p0_y5(45);
	p1_y6(45)<=p0_y6(45);
	p1_y7(45)<=p0_y7(45);
	p1_y8(45)<=p0_y8(45);
	p1_y9(45)<=p0_y9(45);
	p1_y10(45)<=p0_y10(45);
	p1_y0(46)<=p0_y0(46);
	p1_y1(46)<=p0_y1(46);
	p1_y2(46)<=p0_y2(46);
	p1_y3(46)<=p0_y3(46);
	p1_y4(46)<=p0_y4(46);
	p1_y5(46)<=p0_y5(46);
	p1_y6(46)<=p0_y6(46);
	p1_y7(46)<=p0_y7(46);
	p1_y8(46)<=p0_y8(46);
	p1_y9(46)<=p0_y9(46);
	p1_y10(46)<=p0_y10(46);
	p1_y0(47)<=p0_y0(47);
	p1_y1(47)<=p0_y1(47);
	p1_y2(47)<=p0_y2(47);
	p1_y3(47)<=p0_y3(47);
	p1_y4(47)<=p0_y4(47);
	p1_y5(47)<=p0_y5(47);
	p1_y6(47)<=p0_y6(47);
	p1_y7(47)<=p0_y7(47);
	p1_y8(47)<=p0_y8(47);
	p1_y9(47)<=p0_y9(47);
	p1_y0(48)<=p0_y0(48);
	p1_y1(48)<=p0_y1(48);
	p1_y2(48)<=p0_y2(48);
	p1_y3(48)<=p0_y3(48);
	p1_y4(48)<=p0_y4(48);
	p1_y5(48)<=p0_y5(48);
	p1_y6(48)<=p0_y6(48);
	p1_y7(48)<=p0_y7(48);
	p1_y8(48)<=p0_y8(48);
	p1_y9(48)<=p0_y9(48);
	p1_y0(49)<=p0_y0(49);
	p1_y1(49)<=p0_y1(49);
	p1_y2(49)<=p0_y2(49);
	p1_y3(49)<=p0_y3(49);
	p1_y4(49)<=p0_y4(49);
	p1_y5(49)<=p0_y5(49);
	p1_y6(49)<=p0_y6(49);
	p1_y7(49)<=p0_y7(49);
	p1_y8(49)<=p0_y8(49);
	p1_y0(50)<=p0_y0(50);
	p1_y1(50)<=p0_y1(50);
	p1_y2(50)<=p0_y2(50);
	p1_y3(50)<=p0_y3(50);
	p1_y4(50)<=p0_y4(50);
	p1_y5(50)<=p0_y5(50);
	p1_y6(50)<=p0_y6(50);
	p1_y7(50)<=p0_y7(50);
	p1_y8(50)<=p0_y8(50);
	p1_y0(51)<=p0_y0(51);
	p1_y1(51)<=p0_y1(51);
	p1_y2(51)<=p0_y2(51);
	p1_y3(51)<=p0_y3(51);
	p1_y4(51)<=p0_y4(51);
	p1_y5(51)<=p0_y5(51);
	p1_y6(51)<=p0_y6(51);
	p1_y7(51)<=p0_y7(51);
	p1_y0(52)<=p0_y0(52);
	p1_y1(52)<=p0_y1(52);
	p1_y2(52)<=p0_y2(52);
	p1_y3(52)<=p0_y3(52);
	p1_y4(52)<=p0_y4(52);
	p1_y5(52)<=p0_y5(52);
	p1_y6(52)<=p0_y6(52);
	p1_y7(52)<=p0_y7(52);
	p1_y0(53)<=p0_y0(53);
	p1_y1(53)<=p0_y1(53);
	p1_y2(53)<=p0_y2(53);
	p1_y3(53)<=p0_y3(53);
	p1_y4(53)<=p0_y4(53);
	p1_y5(53)<=p0_y5(53);
	p1_y6(53)<=p0_y6(53);
	p1_y0(54)<=p0_y0(54);
	p1_y1(54)<=p0_y1(54);
	p1_y2(54)<=p0_y2(54);
	p1_y3(54)<=p0_y3(54);
	p1_y4(54)<=p0_y4(54);
	p1_y5(54)<=p0_y5(54);
	p1_y6(54)<=p0_y6(54);
	p1_y0(55)<=p0_y0(55);
	p1_y1(55)<=p0_y1(55);
	p1_y2(55)<=p0_y2(55);
	p1_y3(55)<=p0_y3(55);
	p1_y4(55)<=p0_y4(55);
	p1_y5(55)<=p0_y5(55);
	p1_y0(56)<=p0_y0(56);
	p1_y1(56)<=p0_y1(56);
	p1_y2(56)<=p0_y2(56);
	p1_y3(56)<=p0_y3(56);
	p1_y4(56)<=p0_y4(56);
	p1_y5(56)<=p0_y5(56);
	p1_y0(57)<=p0_y0(57);
	p1_y1(57)<=p0_y1(57);
	p1_y2(57)<=p0_y2(57);
	p1_y3(57)<=p0_y3(57);
	p1_y4(57)<=p0_y4(57);
	p1_y0(58)<=p0_y0(58);
	p1_y1(58)<=p0_y1(58);
	p1_y2(58)<=p0_y2(58);
	p1_y3(58)<=p0_y3(58);
	p1_y4(58)<=p0_y4(58);
	p1_y0(59)<=p0_y0(59);
	p1_y1(59)<=p0_y1(59);
	p1_y2(59)<=p0_y2(59);
	p1_y3(59)<=p0_y3(59);
	p1_y0(60)<=p0_y0(60);
	p1_y1(60)<=p0_y1(60);
	p1_y2(60)<=p0_y2(60);
	p1_y3(60)<=p0_y3(60);
	p1_y0(61)<=p0_y0(61);
	p1_y1(61)<=p0_y1(61);
	p1_y2(61)<=p0_y2(61);
	p1_y0(62)<=p0_y0(62);
	p1_y1(62)<=p0_y1(62);
	p1_y2(62)<=p0_y2(62);
	p1_y0(63)<=p0_y0(63);
	p1_y1(63)<=p0_y1(63);
	p2_y0(0)<=p1_y0(0);
	p2_y1(0)<=p1_y1(0);
	p2_y0(1)<=p1_y0(1);
	p2_y1(1)<=p1_y1(1);
	p2_y0(2)<=p1_y0(2);
	p2_y1(2)<=p1_y1(2);
	p2_y2(2)<=p1_y2(2);
	p2_y0(3)<=p1_y0(3);
	p2_y1(3)<=p1_y1(3);
	p2_y2(3)<=p1_y2(3);
	p2_y0(4)<=p1_y0(4);
	p2_y1(4)<=p1_y1(4);
	p2_y2(4)<=p1_y2(4);
	p2_y3(4)<=p1_y3(4);
	p2_y0(5)<=p1_y0(5);
	p2_y1(5)<=p1_y1(5);
	p2_y2(5)<=p1_y2(5);
	p2_y3(5)<=p1_y3(5);
	p2_y0(6)<=p1_y0(6);
	p2_y1(6)<=p1_y1(6);
	p2_y2(6)<=p1_y2(6);
	p2_y3(6)<=p1_y3(6);
	p2_y4(6)<=p1_y4(6);
	p2_y0(7)<=p1_y0(7);
	p2_y1(7)<=p1_y1(7);
	p2_y2(7)<=p1_y2(7);
	p2_y3(7)<=p1_y3(7);
	p2_y4(7)<=p1_y4(7);
	p2_y0(8)<=p1_y0(8);
	p2_y1(8)<=p1_y1(8);
	p2_y2(8)<=p1_y2(8);
	p2_y3(8)<=p1_y3(8);
	p2_y4(8)<=p1_y4(8);
	p2_y5(8)<=p1_y5(8);
	p2_y0(9)<=p1_y0(9);
	p2_y1(9)<=p1_y1(9);
	p2_y2(9)<=p1_y2(9);
	p2_y3(9)<=p1_y3(9);
	p2_y4(9)<=p1_y4(9);
	p2_y5(9)<=p1_y5(9);
	p2_y0(10)<=p1_y0(10);
	p2_y1(10)<=p1_y1(10);
	p2_y2(10)<=p1_y2(10);
	p2_y3(10)<=p1_y3(10);
	p2_y4(10)<=p1_y4(10);
	p2_y5(10)<=p1_y5(10);
	p2_y6(10)<=p1_y6(10);
	p2_y0(11)<=p1_y0(11);
	p2_y1(11)<=p1_y1(11);
	p2_y2(11)<=p1_y2(11);
	p2_y3(11)<=p1_y3(11);
	p2_y4(11)<=p1_y4(11);
	p2_y5(11)<=p1_y5(11);
	p2_y6(11)<=p1_y6(11);
	p2_y0(12)<=p1_y0(12);
	p2_y1(12)<=p1_y1(12);
	p2_y2(12)<=p1_y2(12);
	p2_y3(12)<=p1_y3(12);
	p2_y4(12)<=p1_y4(12);
	p2_y5(12)<=p1_y5(12);
	p2_y6(12)<=p1_y6(12);
	p2_y7(12)<=p1_y7(12);
	p2_y0(13)<=p1_y0(13);
	p2_y1(13)<=p1_y1(13);
	p2_y2(13)<=p1_y2(13);
	p2_y3(13)<=p1_y3(13);
	p2_y4(13)<=p1_y4(13);
	p2_y5(13)<=p1_y5(13);
	p2_y6(13)<=p1_y6(13);
	p2_y7(13)<=p1_y7(13);
	p2_y0(14)<=p1_y0(14);
	p2_y1(14)<=p1_y1(14);
	p2_y2(14)<=p1_y2(14);
	p2_y3(14)<=p1_y3(14);
	p2_y4(14)<=p1_y4(14);
	p2_y5(14)<=p1_y5(14);
	p2_y6(14)<=p1_y6(14);
	p2_y7(14)<=p1_y7(14);
	p2_y8(14)<=p1_y8(14);
	p2_y0(15)<=p1_y0(15);
	p2_y1(15)<=p1_y1(15);
	p2_y2(15)<=p1_y2(15);
	p2_y3(15)<=p1_y3(15);
	p2_y4(15)<=p1_y4(15);
	p2_y5(15)<=p1_y5(15);
	p2_y6(15)<=p1_y6(15);
	p2_y7(15)<=p1_y7(15);
	p2_y8(15)<=p1_y8(15);
	HA8: HA PORT MAP (p1_y0(16),p1_y1(16),p2_y0(16),p2_y0(17));
	p2_y1(16)<=p1_y2(16);
	p2_y2(16)<=p1_y3(16);
	p2_y3(16)<=p1_y4(16);
	p2_y4(16)<=p1_y5(16);
	p2_y5(16)<=p1_y6(16);
	p2_y6(16)<=p1_y7(16);
	p2_y7(16)<=p1_y8(16);
	p2_y8(16)<=p1_y9(16);
	FA44: FA PORT MAP (p1_y0(17),p1_y1(17),p1_y2(17),p2_y1(17),p2_y0(18));
	p2_y2(17)<=p1_y3(17);
	p2_y3(17)<=p1_y4(17);
	p2_y4(17)<=p1_y5(17);
	p2_y5(17)<=p1_y6(17);
	p2_y6(17)<=p1_y7(17);
	p2_y7(17)<=p1_y8(17);
	p2_y8(17)<=p1_y9(17);
	FA45: FA PORT MAP (p1_y0(18),p1_y1(18),p1_y2(18),p2_y1(18),p2_y0(19));
	HA9: HA PORT MAP (p1_y3(18),p1_y4(18),p2_y2(18),p2_y1(19));
	p2_y3(18)<=p1_y5(18);
	p2_y4(18)<=p1_y6(18);
	p2_y5(18)<=p1_y7(18);
	p2_y6(18)<=p1_y8(18);
	p2_y7(18)<=p1_y9(18);
	p2_y8(18)<=p1_y10(18);
	FA46: FA PORT MAP (p1_y0(19),p1_y1(19),p1_y2(19),p2_y2(19),p2_y0(20));
	FA47: FA PORT MAP (p1_y3(19),p1_y4(19),p1_y5(19),p2_y3(19),p2_y1(20));
	p2_y4(19)<=p1_y6(19);
	p2_y5(19)<=p1_y7(19);
	p2_y6(19)<=p1_y8(19);
	p2_y7(19)<=p1_y9(19);
	p2_y8(19)<=p1_y10(19);
	FA48: FA PORT MAP (p1_y0(20),p1_y1(20),p1_y2(20),p2_y2(20),p2_y0(21));
	FA49: FA PORT MAP (p1_y3(20),p1_y4(20),p1_y5(20),p2_y3(20),p2_y1(21));
	HA10: HA PORT MAP (p1_y6(20),p1_y7(20),p2_y4(20),p2_y2(21));
	p2_y5(20)<=p1_y8(20);
	p2_y6(20)<=p1_y9(20);
	p2_y7(20)<=p1_y10(20);
	p2_y8(20)<=p1_y11(20);
	FA50: FA PORT MAP (p1_y0(21),p1_y1(21),p1_y2(21),p2_y3(21),p2_y0(22));
	FA51: FA PORT MAP (p1_y3(21),p1_y4(21),p1_y5(21),p2_y4(21),p2_y1(22));
	FA52: FA PORT MAP (p1_y6(21),p1_y7(21),p1_y8(21),p2_y5(21),p2_y2(22));
	p2_y6(21)<=p1_y9(21);
	p2_y7(21)<=p1_y10(21);
	p2_y8(21)<=p1_y11(21);
	FA53: FA PORT MAP (p1_y0(22),p1_y1(22),p1_y2(22),p2_y3(22),p2_y0(23));
	FA54: FA PORT MAP (p1_y3(22),p1_y4(22),p1_y5(22),p2_y4(22),p2_y1(23));
	FA55: FA PORT MAP (p1_y6(22),p1_y7(22),p1_y8(22),p2_y5(22),p2_y2(23));
	HA11: HA PORT MAP (p1_y9(22),p1_y10(22),p2_y6(22),p2_y3(23));
	p2_y7(22)<=p1_y11(22);
	p2_y8(22)<=p1_y12(22);
	FA56: FA PORT MAP (p1_y0(23),p1_y1(23),p1_y2(23),p2_y4(23),p2_y0(24));
	FA57: FA PORT MAP (p1_y3(23),p1_y4(23),p1_y5(23),p2_y5(23),p2_y1(24));
	FA58: FA PORT MAP (p1_y6(23),p1_y7(23),p1_y8(23),p2_y6(23),p2_y2(24));
	FA59: FA PORT MAP (p1_y9(23),p1_y10(23),p1_y11(23),p2_y7(23),p2_y3(24));
	p2_y8(23)<=p1_y12(23);
	FA60: FA PORT MAP (p1_y0(24),p1_y1(24),p1_y2(24),p2_y4(24),p2_y0(25));
	FA61: FA PORT MAP (p1_y3(24),p1_y4(24),p1_y5(24),p2_y5(24),p2_y1(25));
	FA62: FA PORT MAP (p1_y6(24),p1_y7(24),p1_y8(24),p2_y6(24),p2_y2(25));
	FA63: FA PORT MAP (p1_y9(24),p1_y10(24),p1_y11(24),p2_y7(24),p2_y3(25));
	p2_y8(24)<=p1_y12(24);
	FA64: FA PORT MAP (p1_y0(25),p1_y1(25),p1_y2(25),p2_y4(25),p2_y0(26));
	FA65: FA PORT MAP (p1_y3(25),p1_y4(25),p1_y5(25),p2_y5(25),p2_y1(26));
	FA66: FA PORT MAP (p1_y6(25),p1_y7(25),p1_y8(25),p2_y6(25),p2_y2(26));
	FA67: FA PORT MAP (p1_y9(25),p1_y10(25),p1_y11(25),p2_y7(25),p2_y3(26));
	p2_y8(25)<=p1_y12(25);
	FA68: FA PORT MAP (p1_y0(26),p1_y1(26),p1_y2(26),p2_y4(26),p2_y0(27));
	FA69: FA PORT MAP (p1_y3(26),p1_y4(26),p1_y5(26),p2_y5(26),p2_y1(27));
	FA70: FA PORT MAP (p1_y6(26),p1_y7(26),p1_y8(26),p2_y6(26),p2_y2(27));
	FA71: FA PORT MAP (p1_y9(26),p1_y10(26),p1_y11(26),p2_y7(26),p2_y3(27));
	p2_y8(26)<=p1_y12(26);
	FA72: FA PORT MAP (p1_y0(27),p1_y1(27),p1_y2(27),p2_y4(27),p2_y0(28));
	FA73: FA PORT MAP (p1_y3(27),p1_y4(27),p1_y5(27),p2_y5(27),p2_y1(28));
	FA74: FA PORT MAP (p1_y6(27),p1_y7(27),p1_y8(27),p2_y6(27),p2_y2(28));
	FA75: FA PORT MAP (p1_y9(27),p1_y10(27),p1_y11(27),p2_y7(27),p2_y3(28));
	p2_y8(27)<=p1_y12(27);
	FA76: FA PORT MAP (p1_y0(28),p1_y1(28),p1_y2(28),p2_y4(28),p2_y0(29));
	FA77: FA PORT MAP (p1_y3(28),p1_y4(28),p1_y5(28),p2_y5(28),p2_y1(29));
	FA78: FA PORT MAP (p1_y6(28),p1_y7(28),p1_y8(28),p2_y6(28),p2_y2(29));
	FA79: FA PORT MAP (p1_y9(28),p1_y10(28),p1_y11(28),p2_y7(28),p2_y3(29));
	p2_y8(28)<=p1_y12(28);
	FA80: FA PORT MAP (p1_y0(29),p1_y1(29),p1_y2(29),p2_y4(29),p2_y0(30));
	FA81: FA PORT MAP (p1_y3(29),p1_y4(29),p1_y5(29),p2_y5(29),p2_y1(30));
	FA82: FA PORT MAP (p1_y6(29),p1_y7(29),p1_y8(29),p2_y6(29),p2_y2(30));
	FA83: FA PORT MAP (p1_y9(29),p1_y10(29),p1_y11(29),p2_y7(29),p2_y3(30));
	p2_y8(29)<=p1_y12(29);
	FA84: FA PORT MAP (p1_y0(30),p1_y1(30),p1_y2(30),p2_y4(30),p2_y0(31));
	FA85: FA PORT MAP (p1_y3(30),p1_y4(30),p1_y5(30),p2_y5(30),p2_y1(31));
	FA86: FA PORT MAP (p1_y6(30),p1_y7(30),p1_y8(30),p2_y6(30),p2_y2(31));
	FA87: FA PORT MAP (p1_y9(30),p1_y10(30),p1_y11(30),p2_y7(30),p2_y3(31));
	p2_y8(30)<=p1_y12(30);
	FA88: FA PORT MAP (p1_y0(31),p1_y1(31),p1_y2(31),p2_y4(31),p2_y0(32));
	FA89: FA PORT MAP (p1_y3(31),p1_y4(31),p1_y5(31),p2_y5(31),p2_y1(32));
	FA90: FA PORT MAP (p1_y6(31),p1_y7(31),p1_y8(31),p2_y6(31),p2_y2(32));
	FA91: FA PORT MAP (p1_y9(31),p1_y10(31),p1_y11(31),p2_y7(31),p2_y3(32));
	p2_y8(31)<=p1_y12(31);
	FA92: FA PORT MAP (p1_y0(32),p1_y1(32),p1_y2(32),p2_y4(32),p2_y0(33));
	FA93: FA PORT MAP (p1_y3(32),p1_y4(32),p1_y5(32),p2_y5(32),p2_y1(33));
	FA94: FA PORT MAP (p1_y6(32),p1_y7(32),p1_y8(32),p2_y6(32),p2_y2(33));
	FA95: FA PORT MAP (p1_y9(32),p1_y10(32),p1_y11(32),p2_y7(32),p2_y3(33));
	p2_y8(32)<=p1_y12(32);
	FA96: FA PORT MAP (p1_y0(33),p1_y1(33),p1_y2(33),p2_y4(33),p2_y0(34));
	FA97: FA PORT MAP (p1_y3(33),p1_y4(33),p1_y5(33),p2_y5(33),p2_y1(34));
	FA98: FA PORT MAP (p1_y6(33),p1_y7(33),p1_y8(33),p2_y6(33),p2_y2(34));
	FA99: FA PORT MAP (p1_y9(33),p1_y10(33),p1_y11(33),p2_y7(33),p2_y3(34));
	p2_y8(33)<=p1_y12(33);
	FA100: FA PORT MAP (p1_y0(34),p1_y1(34),p1_y2(34),p2_y4(34),p2_y0(35));
	FA101: FA PORT MAP (p1_y3(34),p1_y4(34),p1_y5(34),p2_y5(34),p2_y1(35));
	FA102: FA PORT MAP (p1_y6(34),p1_y7(34),p1_y8(34),p2_y6(34),p2_y2(35));
	FA103: FA PORT MAP (p1_y9(34),p1_y10(34),p1_y11(34),p2_y7(34),p2_y3(35));
	p2_y8(34)<=p1_y12(34);
	FA104: FA PORT MAP (p1_y0(35),p1_y1(35),p1_y2(35),p2_y4(35),p2_y0(36));
	FA105: FA PORT MAP (p1_y3(35),p1_y4(35),p1_y5(35),p2_y5(35),p2_y1(36));
	FA106: FA PORT MAP (p1_y6(35),p1_y7(35),p1_y8(35),p2_y6(35),p2_y2(36));
	FA107: FA PORT MAP (p1_y9(35),p1_y10(35),p1_y11(35),p2_y7(35),p2_y3(36));
	p2_y8(35)<=p1_y12(35);
	FA108: FA PORT MAP (p1_y0(36),p1_y1(36),p1_y2(36),p2_y4(36),p2_y0(37));
	FA109: FA PORT MAP (p1_y3(36),p1_y4(36),p1_y5(36),p2_y5(36),p2_y1(37));
	FA110: FA PORT MAP (p1_y6(36),p1_y7(36),p1_y8(36),p2_y6(36),p2_y2(37));
	FA111: FA PORT MAP (p1_y9(36),p1_y10(36),p1_y11(36),p2_y7(36),p2_y3(37));
	p2_y8(36)<=p1_y12(36);
	FA112: FA PORT MAP (p1_y0(37),p1_y1(37),p1_y2(37),p2_y4(37),p2_y0(38));
	FA113: FA PORT MAP (p1_y3(37),p1_y4(37),p1_y5(37),p2_y5(37),p2_y1(38));
	FA114: FA PORT MAP (p1_y6(37),p1_y7(37),p1_y8(37),p2_y6(37),p2_y2(38));
	FA115: FA PORT MAP (p1_y9(37),p1_y10(37),p1_y11(37),p2_y7(37),p2_y3(38));
	p2_y8(37)<=p1_y12(37);
	FA116: FA PORT MAP (p1_y0(38),p1_y1(38),p1_y2(38),p2_y4(38),p2_y0(39));
	FA117: FA PORT MAP (p1_y3(38),p1_y4(38),p1_y5(38),p2_y5(38),p2_y1(39));
	FA118: FA PORT MAP (p1_y6(38),p1_y7(38),p1_y8(38),p2_y6(38),p2_y2(39));
	FA119: FA PORT MAP (p1_y9(38),p1_y10(38),p1_y11(38),p2_y7(38),p2_y3(39));
	p2_y8(38)<=p1_y12(38);
	FA120: FA PORT MAP (p1_y0(39),p1_y1(39),p1_y2(39),p2_y4(39),p2_y0(40));
	FA121: FA PORT MAP (p1_y3(39),p1_y4(39),p1_y5(39),p2_y5(39),p2_y1(40));
	FA122: FA PORT MAP (p1_y6(39),p1_y7(39),p1_y8(39),p2_y6(39),p2_y2(40));
	FA123: FA PORT MAP (p1_y9(39),p1_y10(39),p1_y11(39),p2_y7(39),p2_y3(40));
	p2_y8(39)<=p1_y12(39);
	FA124: FA PORT MAP (p1_y0(40),p1_y1(40),p1_y2(40),p2_y4(40),p2_y0(41));
	FA125: FA PORT MAP (p1_y3(40),p1_y4(40),p1_y5(40),p2_y5(40),p2_y1(41));
	FA126: FA PORT MAP (p1_y6(40),p1_y7(40),p1_y8(40),p2_y6(40),p2_y2(41));
	FA127: FA PORT MAP (p1_y9(40),p1_y10(40),p1_y11(40),p2_y7(40),p2_y3(41));
	p2_y8(40)<=p1_y12(40);
	FA128: FA PORT MAP (p1_y0(41),p1_y1(41),p1_y2(41),p2_y4(41),p2_y0(42));
	FA129: FA PORT MAP (p1_y3(41),p1_y4(41),p1_y5(41),p2_y5(41),p2_y1(42));
	FA130: FA PORT MAP (p1_y6(41),p1_y7(41),p1_y8(41),p2_y6(41),p2_y2(42));
	FA131: FA PORT MAP (p1_y9(41),p1_y10(41),p1_y11(41),p2_y7(41),p2_y3(42));
	p2_y8(41)<=p1_y12(41);
	FA132: FA PORT MAP (p1_y0(42),p1_y1(42),p1_y2(42),p2_y4(42),p2_y0(43));
	FA133: FA PORT MAP (p1_y3(42),p1_y4(42),p1_y5(42),p2_y5(42),p2_y1(43));
	FA134: FA PORT MAP (p1_y6(42),p1_y7(42),p1_y8(42),p2_y6(42),p2_y2(43));
	FA135: FA PORT MAP (p1_y9(42),p1_y10(42),p1_y11(42),p2_y7(42),p2_y3(43));
	p2_y8(42)<=p1_y12(42);
	FA136: FA PORT MAP (p1_y0(43),p1_y1(43),p1_y2(43),p2_y4(43),p2_y0(44));
	FA137: FA PORT MAP (p1_y3(43),p1_y4(43),p1_y5(43),p2_y5(43),p2_y1(44));
	FA138: FA PORT MAP (p1_y6(43),p1_y7(43),p1_y8(43),p2_y6(43),p2_y2(44));
	FA139: FA PORT MAP (p1_y9(43),p1_y10(43),p1_y11(43),p2_y7(43),p2_y3(44));
	p2_y8(43)<=p1_y12(43);
	FA140: FA PORT MAP (p1_y0(44),p1_y1(44),p1_y2(44),p2_y4(44),p2_y0(45));
	FA141: FA PORT MAP (p1_y3(44),p1_y4(44),p1_y5(44),p2_y5(44),p2_y1(45));
	FA142: FA PORT MAP (p1_y6(44),p1_y7(44),p1_y8(44),p2_y6(44),p2_y2(45));
	HA12: HA PORT MAP (p1_y9(44),p1_y10(44),p2_y7(44),p2_y3(45));
	p2_y8(44)<=p1_y11(44);
	FA143: FA PORT MAP (p1_y0(45),p1_y1(45),p1_y2(45),p2_y4(45),p2_y0(46));
	FA144: FA PORT MAP (p1_y3(45),p1_y4(45),p1_y5(45),p2_y5(45),p2_y1(46));
	FA145: FA PORT MAP (p1_y6(45),p1_y7(45),p1_y8(45),p2_y6(45),p2_y2(46));
	p2_y7(45)<=p1_y9(45);
	p2_y8(45)<=p1_y10(45);
	FA146: FA PORT MAP (p1_y0(46),p1_y1(46),p1_y2(46),p2_y3(46),p2_y0(47));
	FA147: FA PORT MAP (p1_y3(46),p1_y4(46),p1_y5(46),p2_y4(46),p2_y1(47));
	HA13: HA PORT MAP (p1_y6(46),p1_y7(46),p2_y5(46),p2_y2(47));
	p2_y6(46)<=p1_y8(46);
	p2_y7(46)<=p1_y9(46);
	p2_y8(46)<=p1_y10(46);
	FA148: FA PORT MAP (p1_y0(47),p1_y1(47),p1_y2(47),p2_y3(47),p2_y0(48));
	FA149: FA PORT MAP (p1_y3(47),p1_y4(47),p1_y5(47),p2_y4(47),p2_y1(48));
	p2_y5(47)<=p1_y6(47);
	p2_y6(47)<=p1_y7(47);
	p2_y7(47)<=p1_y8(47);
	p2_y8(47)<=p1_y9(47);
	FA150: FA PORT MAP (p1_y0(48),p1_y1(48),p1_y2(48),p2_y2(48),p2_y0(49));
	HA14: HA PORT MAP (p1_y3(48),p1_y4(48),p2_y3(48),p2_y1(49));
	p2_y4(48)<=p1_y5(48);
	p2_y5(48)<=p1_y6(48);
	p2_y6(48)<=p1_y7(48);
	p2_y7(48)<=p1_y8(48);
	p2_y8(48)<=p1_y9(48);
	FA151: FA PORT MAP (p1_y0(49),p1_y1(49),p1_y2(49),p2_y2(49),p2_y0(50));
	p2_y3(49)<=p1_y3(49);
	p2_y4(49)<=p1_y4(49);
	p2_y5(49)<=p1_y5(49);
	p2_y6(49)<=p1_y6(49);
	p2_y7(49)<=p1_y7(49);
	p2_y8(49)<=p1_y8(49);
	HA15: HA PORT MAP (p1_y0(50),p1_y1(50),p2_y1(50),p2_y0(51));
	p2_y2(50)<=p1_y2(50);
	p2_y3(50)<=p1_y3(50);
	p2_y4(50)<=p1_y4(50);
	p2_y5(50)<=p1_y5(50);
	p2_y6(50)<=p1_y6(50);
	p2_y7(50)<=p1_y7(50);
	p2_y8(50)<=p1_y8(50);
	p2_y1(51)<=p1_y0(51);
	p2_y2(51)<=p1_y1(51);
	p2_y3(51)<=p1_y2(51);
	p2_y4(51)<=p1_y3(51);
	p2_y5(51)<=p1_y4(51);
	p2_y6(51)<=p1_y5(51);
	p2_y7(51)<=p1_y6(51);
	p2_y8(51)<=p1_y7(51);
	p2_y0(52)<=p1_y0(52);
	p2_y1(52)<=p1_y1(52);
	p2_y2(52)<=p1_y2(52);
	p2_y3(52)<=p1_y3(52);
	p2_y4(52)<=p1_y4(52);
	p2_y5(52)<=p1_y5(52);
	p2_y6(52)<=p1_y6(52);
	p2_y7(52)<=p1_y7(52);
	p2_y0(53)<=p1_y0(53);
	p2_y1(53)<=p1_y1(53);
	p2_y2(53)<=p1_y2(53);
	p2_y3(53)<=p1_y3(53);
	p2_y4(53)<=p1_y4(53);
	p2_y5(53)<=p1_y5(53);
	p2_y6(53)<=p1_y6(53);
	p2_y0(54)<=p1_y0(54);
	p2_y1(54)<=p1_y1(54);
	p2_y2(54)<=p1_y2(54);
	p2_y3(54)<=p1_y3(54);
	p2_y4(54)<=p1_y4(54);
	p2_y5(54)<=p1_y5(54);
	p2_y6(54)<=p1_y6(54);
	p2_y0(55)<=p1_y0(55);
	p2_y1(55)<=p1_y1(55);
	p2_y2(55)<=p1_y2(55);
	p2_y3(55)<=p1_y3(55);
	p2_y4(55)<=p1_y4(55);
	p2_y5(55)<=p1_y5(55);
	p2_y0(56)<=p1_y0(56);
	p2_y1(56)<=p1_y1(56);
	p2_y2(56)<=p1_y2(56);
	p2_y3(56)<=p1_y3(56);
	p2_y4(56)<=p1_y4(56);
	p2_y5(56)<=p1_y5(56);
	p2_y0(57)<=p1_y0(57);
	p2_y1(57)<=p1_y1(57);
	p2_y2(57)<=p1_y2(57);
	p2_y3(57)<=p1_y3(57);
	p2_y4(57)<=p1_y4(57);
	p2_y0(58)<=p1_y0(58);
	p2_y1(58)<=p1_y1(58);
	p2_y2(58)<=p1_y2(58);
	p2_y3(58)<=p1_y3(58);
	p2_y4(58)<=p1_y4(58);
	p2_y0(59)<=p1_y0(59);
	p2_y1(59)<=p1_y1(59);
	p2_y2(59)<=p1_y2(59);
	p2_y3(59)<=p1_y3(59);
	p2_y0(60)<=p1_y0(60);
	p2_y1(60)<=p1_y1(60);
	p2_y2(60)<=p1_y2(60);
	p2_y3(60)<=p1_y3(60);
	p2_y0(61)<=p1_y0(61);
	p2_y1(61)<=p1_y1(61);
	p2_y2(61)<=p1_y2(61);
	p2_y0(62)<=p1_y0(62);
	p2_y1(62)<=p1_y1(62);
	p2_y2(62)<=p1_y2(62);
	p2_y0(63)<=p1_y0(63);
	p2_y1(63)<=p1_y1(63);
	p3_y0(0)<=p2_y0(0);
	p3_y1(0)<=p2_y1(0);
	p3_y0(1)<=p2_y0(1);
	p3_y1(1)<=p2_y1(1);
	p3_y0(2)<=p2_y0(2);
	p3_y1(2)<=p2_y1(2);
	p3_y2(2)<=p2_y2(2);
	p3_y0(3)<=p2_y0(3);
	p3_y1(3)<=p2_y1(3);
	p3_y2(3)<=p2_y2(3);
	p3_y0(4)<=p2_y0(4);
	p3_y1(4)<=p2_y1(4);
	p3_y2(4)<=p2_y2(4);
	p3_y3(4)<=p2_y3(4);
	p3_y0(5)<=p2_y0(5);
	p3_y1(5)<=p2_y1(5);
	p3_y2(5)<=p2_y2(5);
	p3_y3(5)<=p2_y3(5);
	p3_y0(6)<=p2_y0(6);
	p3_y1(6)<=p2_y1(6);
	p3_y2(6)<=p2_y2(6);
	p3_y3(6)<=p2_y3(6);
	p3_y4(6)<=p2_y4(6);
	p3_y0(7)<=p2_y0(7);
	p3_y1(7)<=p2_y1(7);
	p3_y2(7)<=p2_y2(7);
	p3_y3(7)<=p2_y3(7);
	p3_y4(7)<=p2_y4(7);
	p3_y0(8)<=p2_y0(8);
	p3_y1(8)<=p2_y1(8);
	p3_y2(8)<=p2_y2(8);
	p3_y3(8)<=p2_y3(8);
	p3_y4(8)<=p2_y4(8);
	p3_y5(8)<=p2_y5(8);
	p3_y0(9)<=p2_y0(9);
	p3_y1(9)<=p2_y1(9);
	p3_y2(9)<=p2_y2(9);
	p3_y3(9)<=p2_y3(9);
	p3_y4(9)<=p2_y4(9);
	p3_y5(9)<=p2_y5(9);
	HA16: HA PORT MAP (p2_y0(10),p2_y1(10),p3_y0(10),p3_y0(11));
	p3_y1(10)<=p2_y2(10);
	p3_y2(10)<=p2_y3(10);
	p3_y3(10)<=p2_y4(10);
	p3_y4(10)<=p2_y5(10);
	p3_y5(10)<=p2_y6(10);
	FA152: FA PORT MAP (p2_y0(11),p2_y1(11),p2_y2(11),p3_y1(11),p3_y0(12));
	p3_y2(11)<=p2_y3(11);
	p3_y3(11)<=p2_y4(11);
	p3_y4(11)<=p2_y5(11);
	p3_y5(11)<=p2_y6(11);
	FA153: FA PORT MAP (p2_y0(12),p2_y1(12),p2_y2(12),p3_y1(12),p3_y0(13));
	HA17: HA PORT MAP (p2_y3(12),p2_y4(12),p3_y2(12),p3_y1(13));
	p3_y3(12)<=p2_y5(12);
	p3_y4(12)<=p2_y6(12);
	p3_y5(12)<=p2_y7(12);
	FA154: FA PORT MAP (p2_y0(13),p2_y1(13),p2_y2(13),p3_y2(13),p3_y0(14));
	FA155: FA PORT MAP (p2_y3(13),p2_y4(13),p2_y5(13),p3_y3(13),p3_y1(14));
	p3_y4(13)<=p2_y6(13);
	p3_y5(13)<=p2_y7(13);
	FA156: FA PORT MAP (p2_y0(14),p2_y1(14),p2_y2(14),p3_y2(14),p3_y0(15));
	FA157: FA PORT MAP (p2_y3(14),p2_y4(14),p2_y5(14),p3_y3(14),p3_y1(15));
	HA18: HA PORT MAP (p2_y6(14),p2_y7(14),p3_y4(14),p3_y2(15));
	p3_y5(14)<=p2_y8(14);
	FA158: FA PORT MAP (p2_y0(15),p2_y1(15),p2_y2(15),p3_y3(15),p3_y0(16));
	FA159: FA PORT MAP (p2_y3(15),p2_y4(15),p2_y5(15),p3_y4(15),p3_y1(16));
	FA160: FA PORT MAP (p2_y6(15),p2_y7(15),p2_y8(15),p3_y5(15),p3_y2(16));
	FA161: FA PORT MAP (p2_y0(16),p2_y1(16),p2_y2(16),p3_y3(16),p3_y0(17));
	FA162: FA PORT MAP (p2_y3(16),p2_y4(16),p2_y5(16),p3_y4(16),p3_y1(17));
	FA163: FA PORT MAP (p2_y6(16),p2_y7(16),p2_y8(16),p3_y5(16),p3_y2(17));
	FA164: FA PORT MAP (p2_y0(17),p2_y1(17),p2_y2(17),p3_y3(17),p3_y0(18));
	FA165: FA PORT MAP (p2_y3(17),p2_y4(17),p2_y5(17),p3_y4(17),p3_y1(18));
	FA166: FA PORT MAP (p2_y6(17),p2_y7(17),p2_y8(17),p3_y5(17),p3_y2(18));
	FA167: FA PORT MAP (p2_y0(18),p2_y1(18),p2_y2(18),p3_y3(18),p3_y0(19));
	FA168: FA PORT MAP (p2_y3(18),p2_y4(18),p2_y5(18),p3_y4(18),p3_y1(19));
	FA169: FA PORT MAP (p2_y6(18),p2_y7(18),p2_y8(18),p3_y5(18),p3_y2(19));
	FA170: FA PORT MAP (p2_y0(19),p2_y1(19),p2_y2(19),p3_y3(19),p3_y0(20));
	FA171: FA PORT MAP (p2_y3(19),p2_y4(19),p2_y5(19),p3_y4(19),p3_y1(20));
	FA172: FA PORT MAP (p2_y6(19),p2_y7(19),p2_y8(19),p3_y5(19),p3_y2(20));
	FA173: FA PORT MAP (p2_y0(20),p2_y1(20),p2_y2(20),p3_y3(20),p3_y0(21));
	FA174: FA PORT MAP (p2_y3(20),p2_y4(20),p2_y5(20),p3_y4(20),p3_y1(21));
	FA175: FA PORT MAP (p2_y6(20),p2_y7(20),p2_y8(20),p3_y5(20),p3_y2(21));
	FA176: FA PORT MAP (p2_y0(21),p2_y1(21),p2_y2(21),p3_y3(21),p3_y0(22));
	FA177: FA PORT MAP (p2_y3(21),p2_y4(21),p2_y5(21),p3_y4(21),p3_y1(22));
	FA178: FA PORT MAP (p2_y6(21),p2_y7(21),p2_y8(21),p3_y5(21),p3_y2(22));
	FA179: FA PORT MAP (p2_y0(22),p2_y1(22),p2_y2(22),p3_y3(22),p3_y0(23));
	FA180: FA PORT MAP (p2_y3(22),p2_y4(22),p2_y5(22),p3_y4(22),p3_y1(23));
	FA181: FA PORT MAP (p2_y6(22),p2_y7(22),p2_y8(22),p3_y5(22),p3_y2(23));
	FA182: FA PORT MAP (p2_y0(23),p2_y1(23),p2_y2(23),p3_y3(23),p3_y0(24));
	FA183: FA PORT MAP (p2_y3(23),p2_y4(23),p2_y5(23),p3_y4(23),p3_y1(24));
	FA184: FA PORT MAP (p2_y6(23),p2_y7(23),p2_y8(23),p3_y5(23),p3_y2(24));
	FA185: FA PORT MAP (p2_y0(24),p2_y1(24),p2_y2(24),p3_y3(24),p3_y0(25));
	FA186: FA PORT MAP (p2_y3(24),p2_y4(24),p2_y5(24),p3_y4(24),p3_y1(25));
	FA187: FA PORT MAP (p2_y6(24),p2_y7(24),p2_y8(24),p3_y5(24),p3_y2(25));
	FA188: FA PORT MAP (p2_y0(25),p2_y1(25),p2_y2(25),p3_y3(25),p3_y0(26));
	FA189: FA PORT MAP (p2_y3(25),p2_y4(25),p2_y5(25),p3_y4(25),p3_y1(26));
	FA190: FA PORT MAP (p2_y6(25),p2_y7(25),p2_y8(25),p3_y5(25),p3_y2(26));
	FA191: FA PORT MAP (p2_y0(26),p2_y1(26),p2_y2(26),p3_y3(26),p3_y0(27));
	FA192: FA PORT MAP (p2_y3(26),p2_y4(26),p2_y5(26),p3_y4(26),p3_y1(27));
	FA193: FA PORT MAP (p2_y6(26),p2_y7(26),p2_y8(26),p3_y5(26),p3_y2(27));
	FA194: FA PORT MAP (p2_y0(27),p2_y1(27),p2_y2(27),p3_y3(27),p3_y0(28));
	FA195: FA PORT MAP (p2_y3(27),p2_y4(27),p2_y5(27),p3_y4(27),p3_y1(28));
	FA196: FA PORT MAP (p2_y6(27),p2_y7(27),p2_y8(27),p3_y5(27),p3_y2(28));
	FA197: FA PORT MAP (p2_y0(28),p2_y1(28),p2_y2(28),p3_y3(28),p3_y0(29));
	FA198: FA PORT MAP (p2_y3(28),p2_y4(28),p2_y5(28),p3_y4(28),p3_y1(29));
	FA199: FA PORT MAP (p2_y6(28),p2_y7(28),p2_y8(28),p3_y5(28),p3_y2(29));
	FA200: FA PORT MAP (p2_y0(29),p2_y1(29),p2_y2(29),p3_y3(29),p3_y0(30));
	FA201: FA PORT MAP (p2_y3(29),p2_y4(29),p2_y5(29),p3_y4(29),p3_y1(30));
	FA202: FA PORT MAP (p2_y6(29),p2_y7(29),p2_y8(29),p3_y5(29),p3_y2(30));
	FA203: FA PORT MAP (p2_y0(30),p2_y1(30),p2_y2(30),p3_y3(30),p3_y0(31));
	FA204: FA PORT MAP (p2_y3(30),p2_y4(30),p2_y5(30),p3_y4(30),p3_y1(31));
	FA205: FA PORT MAP (p2_y6(30),p2_y7(30),p2_y8(30),p3_y5(30),p3_y2(31));
	FA206: FA PORT MAP (p2_y0(31),p2_y1(31),p2_y2(31),p3_y3(31),p3_y0(32));
	FA207: FA PORT MAP (p2_y3(31),p2_y4(31),p2_y5(31),p3_y4(31),p3_y1(32));
	FA208: FA PORT MAP (p2_y6(31),p2_y7(31),p2_y8(31),p3_y5(31),p3_y2(32));
	FA209: FA PORT MAP (p2_y0(32),p2_y1(32),p2_y2(32),p3_y3(32),p3_y0(33));
	FA210: FA PORT MAP (p2_y3(32),p2_y4(32),p2_y5(32),p3_y4(32),p3_y1(33));
	FA211: FA PORT MAP (p2_y6(32),p2_y7(32),p2_y8(32),p3_y5(32),p3_y2(33));
	FA212: FA PORT MAP (p2_y0(33),p2_y1(33),p2_y2(33),p3_y3(33),p3_y0(34));
	FA213: FA PORT MAP (p2_y3(33),p2_y4(33),p2_y5(33),p3_y4(33),p3_y1(34));
	FA214: FA PORT MAP (p2_y6(33),p2_y7(33),p2_y8(33),p3_y5(33),p3_y2(34));
	FA215: FA PORT MAP (p2_y0(34),p2_y1(34),p2_y2(34),p3_y3(34),p3_y0(35));
	FA216: FA PORT MAP (p2_y3(34),p2_y4(34),p2_y5(34),p3_y4(34),p3_y1(35));
	FA217: FA PORT MAP (p2_y6(34),p2_y7(34),p2_y8(34),p3_y5(34),p3_y2(35));
	FA218: FA PORT MAP (p2_y0(35),p2_y1(35),p2_y2(35),p3_y3(35),p3_y0(36));
	FA219: FA PORT MAP (p2_y3(35),p2_y4(35),p2_y5(35),p3_y4(35),p3_y1(36));
	FA220: FA PORT MAP (p2_y6(35),p2_y7(35),p2_y8(35),p3_y5(35),p3_y2(36));
	FA221: FA PORT MAP (p2_y0(36),p2_y1(36),p2_y2(36),p3_y3(36),p3_y0(37));
	FA222: FA PORT MAP (p2_y3(36),p2_y4(36),p2_y5(36),p3_y4(36),p3_y1(37));
	FA223: FA PORT MAP (p2_y6(36),p2_y7(36),p2_y8(36),p3_y5(36),p3_y2(37));
	FA224: FA PORT MAP (p2_y0(37),p2_y1(37),p2_y2(37),p3_y3(37),p3_y0(38));
	FA225: FA PORT MAP (p2_y3(37),p2_y4(37),p2_y5(37),p3_y4(37),p3_y1(38));
	FA226: FA PORT MAP (p2_y6(37),p2_y7(37),p2_y8(37),p3_y5(37),p3_y2(38));
	FA227: FA PORT MAP (p2_y0(38),p2_y1(38),p2_y2(38),p3_y3(38),p3_y0(39));
	FA228: FA PORT MAP (p2_y3(38),p2_y4(38),p2_y5(38),p3_y4(38),p3_y1(39));
	FA229: FA PORT MAP (p2_y6(38),p2_y7(38),p2_y8(38),p3_y5(38),p3_y2(39));
	FA230: FA PORT MAP (p2_y0(39),p2_y1(39),p2_y2(39),p3_y3(39),p3_y0(40));
	FA231: FA PORT MAP (p2_y3(39),p2_y4(39),p2_y5(39),p3_y4(39),p3_y1(40));
	FA232: FA PORT MAP (p2_y6(39),p2_y7(39),p2_y8(39),p3_y5(39),p3_y2(40));
	FA233: FA PORT MAP (p2_y0(40),p2_y1(40),p2_y2(40),p3_y3(40),p3_y0(41));
	FA234: FA PORT MAP (p2_y3(40),p2_y4(40),p2_y5(40),p3_y4(40),p3_y1(41));
	FA235: FA PORT MAP (p2_y6(40),p2_y7(40),p2_y8(40),p3_y5(40),p3_y2(41));
	FA236: FA PORT MAP (p2_y0(41),p2_y1(41),p2_y2(41),p3_y3(41),p3_y0(42));
	FA237: FA PORT MAP (p2_y3(41),p2_y4(41),p2_y5(41),p3_y4(41),p3_y1(42));
	FA238: FA PORT MAP (p2_y6(41),p2_y7(41),p2_y8(41),p3_y5(41),p3_y2(42));
	FA239: FA PORT MAP (p2_y0(42),p2_y1(42),p2_y2(42),p3_y3(42),p3_y0(43));
	FA240: FA PORT MAP (p2_y3(42),p2_y4(42),p2_y5(42),p3_y4(42),p3_y1(43));
	FA241: FA PORT MAP (p2_y6(42),p2_y7(42),p2_y8(42),p3_y5(42),p3_y2(43));
	FA242: FA PORT MAP (p2_y0(43),p2_y1(43),p2_y2(43),p3_y3(43),p3_y0(44));
	FA243: FA PORT MAP (p2_y3(43),p2_y4(43),p2_y5(43),p3_y4(43),p3_y1(44));
	FA244: FA PORT MAP (p2_y6(43),p2_y7(43),p2_y8(43),p3_y5(43),p3_y2(44));
	FA245: FA PORT MAP (p2_y0(44),p2_y1(44),p2_y2(44),p3_y3(44),p3_y0(45));
	FA246: FA PORT MAP (p2_y3(44),p2_y4(44),p2_y5(44),p3_y4(44),p3_y1(45));
	FA247: FA PORT MAP (p2_y6(44),p2_y7(44),p2_y8(44),p3_y5(44),p3_y2(45));
	FA248: FA PORT MAP (p2_y0(45),p2_y1(45),p2_y2(45),p3_y3(45),p3_y0(46));
	FA249: FA PORT MAP (p2_y3(45),p2_y4(45),p2_y5(45),p3_y4(45),p3_y1(46));
	FA250: FA PORT MAP (p2_y6(45),p2_y7(45),p2_y8(45),p3_y5(45),p3_y2(46));
	FA251: FA PORT MAP (p2_y0(46),p2_y1(46),p2_y2(46),p3_y3(46),p3_y0(47));
	FA252: FA PORT MAP (p2_y3(46),p2_y4(46),p2_y5(46),p3_y4(46),p3_y1(47));
	FA253: FA PORT MAP (p2_y6(46),p2_y7(46),p2_y8(46),p3_y5(46),p3_y2(47));
	FA254: FA PORT MAP (p2_y0(47),p2_y1(47),p2_y2(47),p3_y3(47),p3_y0(48));
	FA255: FA PORT MAP (p2_y3(47),p2_y4(47),p2_y5(47),p3_y4(47),p3_y1(48));
	FA256: FA PORT MAP (p2_y6(47),p2_y7(47),p2_y8(47),p3_y5(47),p3_y2(48));
	FA257: FA PORT MAP (p2_y0(48),p2_y1(48),p2_y2(48),p3_y3(48),p3_y0(49));
	FA258: FA PORT MAP (p2_y3(48),p2_y4(48),p2_y5(48),p3_y4(48),p3_y1(49));
	FA259: FA PORT MAP (p2_y6(48),p2_y7(48),p2_y8(48),p3_y5(48),p3_y2(49));
	FA260: FA PORT MAP (p2_y0(49),p2_y1(49),p2_y2(49),p3_y3(49),p3_y0(50));
	FA261: FA PORT MAP (p2_y3(49),p2_y4(49),p2_y5(49),p3_y4(49),p3_y1(50));
	FA262: FA PORT MAP (p2_y6(49),p2_y7(49),p2_y8(49),p3_y5(49),p3_y2(50));
	FA263: FA PORT MAP (p2_y0(50),p2_y1(50),p2_y2(50),p3_y3(50),p3_y0(51));
	FA264: FA PORT MAP (p2_y3(50),p2_y4(50),p2_y5(50),p3_y4(50),p3_y1(51));
	FA265: FA PORT MAP (p2_y6(50),p2_y7(50),p2_y8(50),p3_y5(50),p3_y2(51));
	FA266: FA PORT MAP (p2_y0(51),p2_y1(51),p2_y2(51),p3_y3(51),p3_y0(52));
	FA267: FA PORT MAP (p2_y3(51),p2_y4(51),p2_y5(51),p3_y4(51),p3_y1(52));
	FA268: FA PORT MAP (p2_y6(51),p2_y7(51),p2_y8(51),p3_y5(51),p3_y2(52));
	FA269: FA PORT MAP (p2_y0(52),p2_y1(52),p2_y2(52),p3_y3(52),p3_y0(53));
	FA270: FA PORT MAP (p2_y3(52),p2_y4(52),p2_y5(52),p3_y4(52),p3_y1(53));
	HA19: HA PORT MAP (p2_y6(52),p2_y7(52),p3_y5(52),p3_y2(53));
	FA271: FA PORT MAP (p2_y0(53),p2_y1(53),p2_y2(53),p3_y3(53),p3_y0(54));
	FA272: FA PORT MAP (p2_y3(53),p2_y4(53),p2_y5(53),p3_y4(53),p3_y1(54));
	p3_y5(53)<=p2_y6(53);
	FA273: FA PORT MAP (p2_y0(54),p2_y1(54),p2_y2(54),p3_y2(54),p3_y0(55));
	HA20: HA PORT MAP (p2_y3(54),p2_y4(54),p3_y3(54),p3_y1(55));
	p3_y4(54)<=p2_y5(54);
	p3_y5(54)<=p2_y6(54);
	FA274: FA PORT MAP (p2_y0(55),p2_y1(55),p2_y2(55),p3_y2(55),p3_y0(56));
	p3_y3(55)<=p2_y3(55);
	p3_y4(55)<=p2_y4(55);
	p3_y5(55)<=p2_y5(55);
	HA21: HA PORT MAP (p2_y0(56),p2_y1(56),p3_y1(56),p3_y0(57));
	p3_y2(56)<=p2_y2(56);
	p3_y3(56)<=p2_y3(56);
	p3_y4(56)<=p2_y4(56);
	p3_y5(56)<=p2_y5(56);
	p3_y1(57)<=p2_y0(57);
	p3_y2(57)<=p2_y1(57);
	p3_y3(57)<=p2_y2(57);
	p3_y4(57)<=p2_y3(57);
	p3_y5(57)<=p2_y4(57);
	p3_y0(58)<=p2_y0(58);
	p3_y1(58)<=p2_y1(58);
	p3_y2(58)<=p2_y2(58);
	p3_y3(58)<=p2_y3(58);
	p3_y4(58)<=p2_y4(58);
	p3_y0(59)<=p2_y0(59);
	p3_y1(59)<=p2_y1(59);
	p3_y2(59)<=p2_y2(59);
	p3_y3(59)<=p2_y3(59);
	p3_y0(60)<=p2_y0(60);
	p3_y1(60)<=p2_y1(60);
	p3_y2(60)<=p2_y2(60);
	p3_y3(60)<=p2_y3(60);
	p3_y0(61)<=p2_y0(61);
	p3_y1(61)<=p2_y1(61);
	p3_y2(61)<=p2_y2(61);
	p3_y0(62)<=p2_y0(62);
	p3_y1(62)<=p2_y1(62);
	p3_y2(62)<=p2_y2(62);
	p3_y0(63)<=p2_y0(63);
	p3_y1(63)<=p2_y1(63);
	p4_y0(0)<=p3_y0(0);
	p4_y1(0)<=p3_y1(0);
	p4_y0(1)<=p3_y0(1);
	p4_y1(1)<=p3_y1(1);
	p4_y0(2)<=p3_y0(2);
	p4_y1(2)<=p3_y1(2);
	p4_y2(2)<=p3_y2(2);
	p4_y0(3)<=p3_y0(3);
	p4_y1(3)<=p3_y1(3);
	p4_y2(3)<=p3_y2(3);
	p4_y0(4)<=p3_y0(4);
	p4_y1(4)<=p3_y1(4);
	p4_y2(4)<=p3_y2(4);
	p4_y3(4)<=p3_y3(4);
	p4_y0(5)<=p3_y0(5);
	p4_y1(5)<=p3_y1(5);
	p4_y2(5)<=p3_y2(5);
	p4_y3(5)<=p3_y3(5);
	HA22: HA PORT MAP (p3_y0(6),p3_y1(6),p4_y0(6),p4_y0(7));
	p4_y1(6)<=p3_y2(6);
	p4_y2(6)<=p3_y3(6);
	p4_y3(6)<=p3_y4(6);
	FA275: FA PORT MAP (p3_y0(7),p3_y1(7),p3_y2(7),p4_y1(7),p4_y0(8));
	p4_y2(7)<=p3_y3(7);
	p4_y3(7)<=p3_y4(7);
	FA276: FA PORT MAP (p3_y0(8),p3_y1(8),p3_y2(8),p4_y1(8),p4_y0(9));
	HA23: HA PORT MAP (p3_y3(8),p3_y4(8),p4_y2(8),p4_y1(9));
	p4_y3(8)<=p3_y5(8);
	FA277: FA PORT MAP (p3_y0(9),p3_y1(9),p3_y2(9),p4_y2(9),p4_y0(10));
	FA278: FA PORT MAP (p3_y3(9),p3_y4(9),p3_y5(9),p4_y3(9),p4_y1(10));
	FA279: FA PORT MAP (p3_y0(10),p3_y1(10),p3_y2(10),p4_y2(10),p4_y0(11));
	FA280: FA PORT MAP (p3_y3(10),p3_y4(10),p3_y5(10),p4_y3(10),p4_y1(11));
	FA281: FA PORT MAP (p3_y0(11),p3_y1(11),p3_y2(11),p4_y2(11),p4_y0(12));
	FA282: FA PORT MAP (p3_y3(11),p3_y4(11),p3_y5(11),p4_y3(11),p4_y1(12));
	FA283: FA PORT MAP (p3_y0(12),p3_y1(12),p3_y2(12),p4_y2(12),p4_y0(13));
	FA284: FA PORT MAP (p3_y3(12),p3_y4(12),p3_y5(12),p4_y3(12),p4_y1(13));
	FA285: FA PORT MAP (p3_y0(13),p3_y1(13),p3_y2(13),p4_y2(13),p4_y0(14));
	FA286: FA PORT MAP (p3_y3(13),p3_y4(13),p3_y5(13),p4_y3(13),p4_y1(14));
	FA287: FA PORT MAP (p3_y0(14),p3_y1(14),p3_y2(14),p4_y2(14),p4_y0(15));
	FA288: FA PORT MAP (p3_y3(14),p3_y4(14),p3_y5(14),p4_y3(14),p4_y1(15));
	FA289: FA PORT MAP (p3_y0(15),p3_y1(15),p3_y2(15),p4_y2(15),p4_y0(16));
	FA290: FA PORT MAP (p3_y3(15),p3_y4(15),p3_y5(15),p4_y3(15),p4_y1(16));
	FA291: FA PORT MAP (p3_y0(16),p3_y1(16),p3_y2(16),p4_y2(16),p4_y0(17));
	FA292: FA PORT MAP (p3_y3(16),p3_y4(16),p3_y5(16),p4_y3(16),p4_y1(17));
	FA293: FA PORT MAP (p3_y0(17),p3_y1(17),p3_y2(17),p4_y2(17),p4_y0(18));
	FA294: FA PORT MAP (p3_y3(17),p3_y4(17),p3_y5(17),p4_y3(17),p4_y1(18));
	FA295: FA PORT MAP (p3_y0(18),p3_y1(18),p3_y2(18),p4_y2(18),p4_y0(19));
	FA296: FA PORT MAP (p3_y3(18),p3_y4(18),p3_y5(18),p4_y3(18),p4_y1(19));
	FA297: FA PORT MAP (p3_y0(19),p3_y1(19),p3_y2(19),p4_y2(19),p4_y0(20));
	FA298: FA PORT MAP (p3_y3(19),p3_y4(19),p3_y5(19),p4_y3(19),p4_y1(20));
	FA299: FA PORT MAP (p3_y0(20),p3_y1(20),p3_y2(20),p4_y2(20),p4_y0(21));
	FA300: FA PORT MAP (p3_y3(20),p3_y4(20),p3_y5(20),p4_y3(20),p4_y1(21));
	FA301: FA PORT MAP (p3_y0(21),p3_y1(21),p3_y2(21),p4_y2(21),p4_y0(22));
	FA302: FA PORT MAP (p3_y3(21),p3_y4(21),p3_y5(21),p4_y3(21),p4_y1(22));
	FA303: FA PORT MAP (p3_y0(22),p3_y1(22),p3_y2(22),p4_y2(22),p4_y0(23));
	FA304: FA PORT MAP (p3_y3(22),p3_y4(22),p3_y5(22),p4_y3(22),p4_y1(23));
	FA305: FA PORT MAP (p3_y0(23),p3_y1(23),p3_y2(23),p4_y2(23),p4_y0(24));
	FA306: FA PORT MAP (p3_y3(23),p3_y4(23),p3_y5(23),p4_y3(23),p4_y1(24));
	FA307: FA PORT MAP (p3_y0(24),p3_y1(24),p3_y2(24),p4_y2(24),p4_y0(25));
	FA308: FA PORT MAP (p3_y3(24),p3_y4(24),p3_y5(24),p4_y3(24),p4_y1(25));
	FA309: FA PORT MAP (p3_y0(25),p3_y1(25),p3_y2(25),p4_y2(25),p4_y0(26));
	FA310: FA PORT MAP (p3_y3(25),p3_y4(25),p3_y5(25),p4_y3(25),p4_y1(26));
	FA311: FA PORT MAP (p3_y0(26),p3_y1(26),p3_y2(26),p4_y2(26),p4_y0(27));
	FA312: FA PORT MAP (p3_y3(26),p3_y4(26),p3_y5(26),p4_y3(26),p4_y1(27));
	FA313: FA PORT MAP (p3_y0(27),p3_y1(27),p3_y2(27),p4_y2(27),p4_y0(28));
	FA314: FA PORT MAP (p3_y3(27),p3_y4(27),p3_y5(27),p4_y3(27),p4_y1(28));
	FA315: FA PORT MAP (p3_y0(28),p3_y1(28),p3_y2(28),p4_y2(28),p4_y0(29));
	FA316: FA PORT MAP (p3_y3(28),p3_y4(28),p3_y5(28),p4_y3(28),p4_y1(29));
	FA317: FA PORT MAP (p3_y0(29),p3_y1(29),p3_y2(29),p4_y2(29),p4_y0(30));
	FA318: FA PORT MAP (p3_y3(29),p3_y4(29),p3_y5(29),p4_y3(29),p4_y1(30));
	FA319: FA PORT MAP (p3_y0(30),p3_y1(30),p3_y2(30),p4_y2(30),p4_y0(31));
	FA320: FA PORT MAP (p3_y3(30),p3_y4(30),p3_y5(30),p4_y3(30),p4_y1(31));
	FA321: FA PORT MAP (p3_y0(31),p3_y1(31),p3_y2(31),p4_y2(31),p4_y0(32));
	FA322: FA PORT MAP (p3_y3(31),p3_y4(31),p3_y5(31),p4_y3(31),p4_y1(32));
	FA323: FA PORT MAP (p3_y0(32),p3_y1(32),p3_y2(32),p4_y2(32),p4_y0(33));
	FA324: FA PORT MAP (p3_y3(32),p3_y4(32),p3_y5(32),p4_y3(32),p4_y1(33));
	FA325: FA PORT MAP (p3_y0(33),p3_y1(33),p3_y2(33),p4_y2(33),p4_y0(34));
	FA326: FA PORT MAP (p3_y3(33),p3_y4(33),p3_y5(33),p4_y3(33),p4_y1(34));
	FA327: FA PORT MAP (p3_y0(34),p3_y1(34),p3_y2(34),p4_y2(34),p4_y0(35));
	FA328: FA PORT MAP (p3_y3(34),p3_y4(34),p3_y5(34),p4_y3(34),p4_y1(35));
	FA329: FA PORT MAP (p3_y0(35),p3_y1(35),p3_y2(35),p4_y2(35),p4_y0(36));
	FA330: FA PORT MAP (p3_y3(35),p3_y4(35),p3_y5(35),p4_y3(35),p4_y1(36));
	FA331: FA PORT MAP (p3_y0(36),p3_y1(36),p3_y2(36),p4_y2(36),p4_y0(37));
	FA332: FA PORT MAP (p3_y3(36),p3_y4(36),p3_y5(36),p4_y3(36),p4_y1(37));
	FA333: FA PORT MAP (p3_y0(37),p3_y1(37),p3_y2(37),p4_y2(37),p4_y0(38));
	FA334: FA PORT MAP (p3_y3(37),p3_y4(37),p3_y5(37),p4_y3(37),p4_y1(38));
	FA335: FA PORT MAP (p3_y0(38),p3_y1(38),p3_y2(38),p4_y2(38),p4_y0(39));
	FA336: FA PORT MAP (p3_y3(38),p3_y4(38),p3_y5(38),p4_y3(38),p4_y1(39));
	FA337: FA PORT MAP (p3_y0(39),p3_y1(39),p3_y2(39),p4_y2(39),p4_y0(40));
	FA338: FA PORT MAP (p3_y3(39),p3_y4(39),p3_y5(39),p4_y3(39),p4_y1(40));
	FA339: FA PORT MAP (p3_y0(40),p3_y1(40),p3_y2(40),p4_y2(40),p4_y0(41));
	FA340: FA PORT MAP (p3_y3(40),p3_y4(40),p3_y5(40),p4_y3(40),p4_y1(41));
	FA341: FA PORT MAP (p3_y0(41),p3_y1(41),p3_y2(41),p4_y2(41),p4_y0(42));
	FA342: FA PORT MAP (p3_y3(41),p3_y4(41),p3_y5(41),p4_y3(41),p4_y1(42));
	FA343: FA PORT MAP (p3_y0(42),p3_y1(42),p3_y2(42),p4_y2(42),p4_y0(43));
	FA344: FA PORT MAP (p3_y3(42),p3_y4(42),p3_y5(42),p4_y3(42),p4_y1(43));
	FA345: FA PORT MAP (p3_y0(43),p3_y1(43),p3_y2(43),p4_y2(43),p4_y0(44));
	FA346: FA PORT MAP (p3_y3(43),p3_y4(43),p3_y5(43),p4_y3(43),p4_y1(44));
	FA347: FA PORT MAP (p3_y0(44),p3_y1(44),p3_y2(44),p4_y2(44),p4_y0(45));
	FA348: FA PORT MAP (p3_y3(44),p3_y4(44),p3_y5(44),p4_y3(44),p4_y1(45));
	FA349: FA PORT MAP (p3_y0(45),p3_y1(45),p3_y2(45),p4_y2(45),p4_y0(46));
	FA350: FA PORT MAP (p3_y3(45),p3_y4(45),p3_y5(45),p4_y3(45),p4_y1(46));
	FA351: FA PORT MAP (p3_y0(46),p3_y1(46),p3_y2(46),p4_y2(46),p4_y0(47));
	FA352: FA PORT MAP (p3_y3(46),p3_y4(46),p3_y5(46),p4_y3(46),p4_y1(47));
	FA353: FA PORT MAP (p3_y0(47),p3_y1(47),p3_y2(47),p4_y2(47),p4_y0(48));
	FA354: FA PORT MAP (p3_y3(47),p3_y4(47),p3_y5(47),p4_y3(47),p4_y1(48));
	FA355: FA PORT MAP (p3_y0(48),p3_y1(48),p3_y2(48),p4_y2(48),p4_y0(49));
	FA356: FA PORT MAP (p3_y3(48),p3_y4(48),p3_y5(48),p4_y3(48),p4_y1(49));
	FA357: FA PORT MAP (p3_y0(49),p3_y1(49),p3_y2(49),p4_y2(49),p4_y0(50));
	FA358: FA PORT MAP (p3_y3(49),p3_y4(49),p3_y5(49),p4_y3(49),p4_y1(50));
	FA359: FA PORT MAP (p3_y0(50),p3_y1(50),p3_y2(50),p4_y2(50),p4_y0(51));
	FA360: FA PORT MAP (p3_y3(50),p3_y4(50),p3_y5(50),p4_y3(50),p4_y1(51));
	FA361: FA PORT MAP (p3_y0(51),p3_y1(51),p3_y2(51),p4_y2(51),p4_y0(52));
	FA362: FA PORT MAP (p3_y3(51),p3_y4(51),p3_y5(51),p4_y3(51),p4_y1(52));
	FA363: FA PORT MAP (p3_y0(52),p3_y1(52),p3_y2(52),p4_y2(52),p4_y0(53));
	FA364: FA PORT MAP (p3_y3(52),p3_y4(52),p3_y5(52),p4_y3(52),p4_y1(53));
	FA365: FA PORT MAP (p3_y0(53),p3_y1(53),p3_y2(53),p4_y2(53),p4_y0(54));
	FA366: FA PORT MAP (p3_y3(53),p3_y4(53),p3_y5(53),p4_y3(53),p4_y1(54));
	FA367: FA PORT MAP (p3_y0(54),p3_y1(54),p3_y2(54),p4_y2(54),p4_y0(55));
	FA368: FA PORT MAP (p3_y3(54),p3_y4(54),p3_y5(54),p4_y3(54),p4_y1(55));
	FA369: FA PORT MAP (p3_y0(55),p3_y1(55),p3_y2(55),p4_y2(55),p4_y0(56));
	FA370: FA PORT MAP (p3_y3(55),p3_y4(55),p3_y5(55),p4_y3(55),p4_y1(56));
	FA371: FA PORT MAP (p3_y0(56),p3_y1(56),p3_y2(56),p4_y2(56),p4_y0(57));
	FA372: FA PORT MAP (p3_y3(56),p3_y4(56),p3_y5(56),p4_y3(56),p4_y1(57));
	FA373: FA PORT MAP (p3_y0(57),p3_y1(57),p3_y2(57),p4_y2(57),p4_y0(58));
	FA374: FA PORT MAP (p3_y3(57),p3_y4(57),p3_y5(57),p4_y3(57),p4_y1(58));
	FA375: FA PORT MAP (p3_y0(58),p3_y1(58),p3_y2(58),p4_y2(58),p4_y0(59));
	HA24: HA PORT MAP (p3_y3(58),p3_y4(58),p4_y3(58),p4_y1(59));
	FA376: FA PORT MAP (p3_y0(59),p3_y1(59),p3_y2(59),p4_y2(59),p4_y0(60));
	p4_y3(59)<=p3_y3(59);
	HA25: HA PORT MAP (p3_y0(60),p3_y1(60),p4_y1(60),p4_y0(61));
	p4_y2(60)<=p3_y2(60);
	p4_y3(60)<=p3_y3(60);
	p4_y1(61)<=p3_y0(61);
	p4_y2(61)<=p3_y1(61);
	p4_y3(61)<=p3_y2(61);
	p4_y0(62)<=p3_y0(62);
	p4_y1(62)<=p3_y1(62);
	p4_y2(62)<=p3_y2(62);
	p4_y0(63)<=p3_y0(63);
	p4_y1(63)<=p3_y1(63);
	p5_y0(0)<=p4_y0(0);
	p5_y1(0)<=p4_y1(0);
	p5_y0(1)<=p4_y0(1);
	p5_y1(1)<=p4_y1(1);
	p5_y0(2)<=p4_y0(2);
	p5_y1(2)<=p4_y1(2);
	p5_y2(2)<=p4_y2(2);
	p5_y0(3)<=p4_y0(3);
	p5_y1(3)<=p4_y1(3);
	p5_y2(3)<=p4_y2(3);
	HA26: HA PORT MAP (p4_y0(4),p4_y1(4),p5_y0(4),p5_y0(5));
	p5_y1(4)<=p4_y2(4);
	p5_y2(4)<=p4_y3(4);
	FA377: FA PORT MAP (p4_y0(5),p4_y1(5),p4_y2(5),p5_y1(5),p5_y0(6));
	p5_y2(5)<=p4_y3(5);
	FA378: FA PORT MAP (p4_y0(6),p4_y1(6),p4_y2(6),p5_y1(6),p5_y0(7));
	p5_y2(6)<=p4_y3(6);
	FA379: FA PORT MAP (p4_y0(7),p4_y1(7),p4_y2(7),p5_y1(7),p5_y0(8));
	p5_y2(7)<=p4_y3(7);
	FA380: FA PORT MAP (p4_y0(8),p4_y1(8),p4_y2(8),p5_y1(8),p5_y0(9));
	p5_y2(8)<=p4_y3(8);
	FA381: FA PORT MAP (p4_y0(9),p4_y1(9),p4_y2(9),p5_y1(9),p5_y0(10));
	p5_y2(9)<=p4_y3(9);
	FA382: FA PORT MAP (p4_y0(10),p4_y1(10),p4_y2(10),p5_y1(10),p5_y0(11));
	p5_y2(10)<=p4_y3(10);
	FA383: FA PORT MAP (p4_y0(11),p4_y1(11),p4_y2(11),p5_y1(11),p5_y0(12));
	p5_y2(11)<=p4_y3(11);
	FA384: FA PORT MAP (p4_y0(12),p4_y1(12),p4_y2(12),p5_y1(12),p5_y0(13));
	p5_y2(12)<=p4_y3(12);
	FA385: FA PORT MAP (p4_y0(13),p4_y1(13),p4_y2(13),p5_y1(13),p5_y0(14));
	p5_y2(13)<=p4_y3(13);
	FA386: FA PORT MAP (p4_y0(14),p4_y1(14),p4_y2(14),p5_y1(14),p5_y0(15));
	p5_y2(14)<=p4_y3(14);
	FA387: FA PORT MAP (p4_y0(15),p4_y1(15),p4_y2(15),p5_y1(15),p5_y0(16));
	p5_y2(15)<=p4_y3(15);
	FA388: FA PORT MAP (p4_y0(16),p4_y1(16),p4_y2(16),p5_y1(16),p5_y0(17));
	p5_y2(16)<=p4_y3(16);
	FA389: FA PORT MAP (p4_y0(17),p4_y1(17),p4_y2(17),p5_y1(17),p5_y0(18));
	p5_y2(17)<=p4_y3(17);
	FA390: FA PORT MAP (p4_y0(18),p4_y1(18),p4_y2(18),p5_y1(18),p5_y0(19));
	p5_y2(18)<=p4_y3(18);
	FA391: FA PORT MAP (p4_y0(19),p4_y1(19),p4_y2(19),p5_y1(19),p5_y0(20));
	p5_y2(19)<=p4_y3(19);
	FA392: FA PORT MAP (p4_y0(20),p4_y1(20),p4_y2(20),p5_y1(20),p5_y0(21));
	p5_y2(20)<=p4_y3(20);
	FA393: FA PORT MAP (p4_y0(21),p4_y1(21),p4_y2(21),p5_y1(21),p5_y0(22));
	p5_y2(21)<=p4_y3(21);
	FA394: FA PORT MAP (p4_y0(22),p4_y1(22),p4_y2(22),p5_y1(22),p5_y0(23));
	p5_y2(22)<=p4_y3(22);
	FA395: FA PORT MAP (p4_y0(23),p4_y1(23),p4_y2(23),p5_y1(23),p5_y0(24));
	p5_y2(23)<=p4_y3(23);
	FA396: FA PORT MAP (p4_y0(24),p4_y1(24),p4_y2(24),p5_y1(24),p5_y0(25));
	p5_y2(24)<=p4_y3(24);
	FA397: FA PORT MAP (p4_y0(25),p4_y1(25),p4_y2(25),p5_y1(25),p5_y0(26));
	p5_y2(25)<=p4_y3(25);
	FA398: FA PORT MAP (p4_y0(26),p4_y1(26),p4_y2(26),p5_y1(26),p5_y0(27));
	p5_y2(26)<=p4_y3(26);
	FA399: FA PORT MAP (p4_y0(27),p4_y1(27),p4_y2(27),p5_y1(27),p5_y0(28));
	p5_y2(27)<=p4_y3(27);
	FA400: FA PORT MAP (p4_y0(28),p4_y1(28),p4_y2(28),p5_y1(28),p5_y0(29));
	p5_y2(28)<=p4_y3(28);
	FA401: FA PORT MAP (p4_y0(29),p4_y1(29),p4_y2(29),p5_y1(29),p5_y0(30));
	p5_y2(29)<=p4_y3(29);
	FA402: FA PORT MAP (p4_y0(30),p4_y1(30),p4_y2(30),p5_y1(30),p5_y0(31));
	p5_y2(30)<=p4_y3(30);
	FA403: FA PORT MAP (p4_y0(31),p4_y1(31),p4_y2(31),p5_y1(31),p5_y0(32));
	p5_y2(31)<=p4_y3(31);
	FA404: FA PORT MAP (p4_y0(32),p4_y1(32),p4_y2(32),p5_y1(32),p5_y0(33));
	p5_y2(32)<=p4_y3(32);
	FA405: FA PORT MAP (p4_y0(33),p4_y1(33),p4_y2(33),p5_y1(33),p5_y0(34));
	p5_y2(33)<=p4_y3(33);
	FA406: FA PORT MAP (p4_y0(34),p4_y1(34),p4_y2(34),p5_y1(34),p5_y0(35));
	p5_y2(34)<=p4_y3(34);
	FA407: FA PORT MAP (p4_y0(35),p4_y1(35),p4_y2(35),p5_y1(35),p5_y0(36));
	p5_y2(35)<=p4_y3(35);
	FA408: FA PORT MAP (p4_y0(36),p4_y1(36),p4_y2(36),p5_y1(36),p5_y0(37));
	p5_y2(36)<=p4_y3(36);
	FA409: FA PORT MAP (p4_y0(37),p4_y1(37),p4_y2(37),p5_y1(37),p5_y0(38));
	p5_y2(37)<=p4_y3(37);
	FA410: FA PORT MAP (p4_y0(38),p4_y1(38),p4_y2(38),p5_y1(38),p5_y0(39));
	p5_y2(38)<=p4_y3(38);
	FA411: FA PORT MAP (p4_y0(39),p4_y1(39),p4_y2(39),p5_y1(39),p5_y0(40));
	p5_y2(39)<=p4_y3(39);
	FA412: FA PORT MAP (p4_y0(40),p4_y1(40),p4_y2(40),p5_y1(40),p5_y0(41));
	p5_y2(40)<=p4_y3(40);
	FA413: FA PORT MAP (p4_y0(41),p4_y1(41),p4_y2(41),p5_y1(41),p5_y0(42));
	p5_y2(41)<=p4_y3(41);
	FA414: FA PORT MAP (p4_y0(42),p4_y1(42),p4_y2(42),p5_y1(42),p5_y0(43));
	p5_y2(42)<=p4_y3(42);
	FA415: FA PORT MAP (p4_y0(43),p4_y1(43),p4_y2(43),p5_y1(43),p5_y0(44));
	p5_y2(43)<=p4_y3(43);
	FA416: FA PORT MAP (p4_y0(44),p4_y1(44),p4_y2(44),p5_y1(44),p5_y0(45));
	p5_y2(44)<=p4_y3(44);
	FA417: FA PORT MAP (p4_y0(45),p4_y1(45),p4_y2(45),p5_y1(45),p5_y0(46));
	p5_y2(45)<=p4_y3(45);
	FA418: FA PORT MAP (p4_y0(46),p4_y1(46),p4_y2(46),p5_y1(46),p5_y0(47));
	p5_y2(46)<=p4_y3(46);
	FA419: FA PORT MAP (p4_y0(47),p4_y1(47),p4_y2(47),p5_y1(47),p5_y0(48));
	p5_y2(47)<=p4_y3(47);
	FA420: FA PORT MAP (p4_y0(48),p4_y1(48),p4_y2(48),p5_y1(48),p5_y0(49));
	p5_y2(48)<=p4_y3(48);
	FA421: FA PORT MAP (p4_y0(49),p4_y1(49),p4_y2(49),p5_y1(49),p5_y0(50));
	p5_y2(49)<=p4_y3(49);
	FA422: FA PORT MAP (p4_y0(50),p4_y1(50),p4_y2(50),p5_y1(50),p5_y0(51));
	p5_y2(50)<=p4_y3(50);
	FA423: FA PORT MAP (p4_y0(51),p4_y1(51),p4_y2(51),p5_y1(51),p5_y0(52));
	p5_y2(51)<=p4_y3(51);
	FA424: FA PORT MAP (p4_y0(52),p4_y1(52),p4_y2(52),p5_y1(52),p5_y0(53));
	p5_y2(52)<=p4_y3(52);
	FA425: FA PORT MAP (p4_y0(53),p4_y1(53),p4_y2(53),p5_y1(53),p5_y0(54));
	p5_y2(53)<=p4_y3(53);
	FA426: FA PORT MAP (p4_y0(54),p4_y1(54),p4_y2(54),p5_y1(54),p5_y0(55));
	p5_y2(54)<=p4_y3(54);
	FA427: FA PORT MAP (p4_y0(55),p4_y1(55),p4_y2(55),p5_y1(55),p5_y0(56));
	p5_y2(55)<=p4_y3(55);
	FA428: FA PORT MAP (p4_y0(56),p4_y1(56),p4_y2(56),p5_y1(56),p5_y0(57));
	p5_y2(56)<=p4_y3(56);
	FA429: FA PORT MAP (p4_y0(57),p4_y1(57),p4_y2(57),p5_y1(57),p5_y0(58));
	p5_y2(57)<=p4_y3(57);
	FA430: FA PORT MAP (p4_y0(58),p4_y1(58),p4_y2(58),p5_y1(58),p5_y0(59));
	p5_y2(58)<=p4_y3(58);
	FA431: FA PORT MAP (p4_y0(59),p4_y1(59),p4_y2(59),p5_y1(59),p5_y0(60));
	p5_y2(59)<=p4_y3(59);
	FA432: FA PORT MAP (p4_y0(60),p4_y1(60),p4_y2(60),p5_y1(60),p5_y0(61));
	p5_y2(60)<=p4_y3(60);
	FA433: FA PORT MAP (p4_y0(61),p4_y1(61),p4_y2(61),p5_y1(61),p5_y0(62));
	p5_y2(61)<=p4_y3(61);
	HA27: HA PORT MAP (p4_y0(62),p4_y1(62),p5_y1(62),p5_y0(63));
	p5_y2(62)<=p4_y2(62);
	p5_y1(63)<=p4_y0(63);
	p5_y2(63)<=p4_y1(63);
	p6_y0(0)<=p5_y0(0);
	p6_y1(0)<=p5_y1(0);
	p6_y0(1)<=p5_y0(1);
	p6_y1(1)<=p5_y1(1);
	HA28: HA PORT MAP (p5_y0(2),p5_y1(2),p6_y0(2),p6_y0(3));
	p6_y1(2)<=p5_y2(2);
	FA434: FA PORT MAP (p5_y0(3),p5_y1(3),p5_y2(3),p6_y1(3),p6_y0(4));
	FA435: FA PORT MAP (p5_y0(4),p5_y1(4),p5_y2(4),p6_y1(4),p6_y0(5));
	FA436: FA PORT MAP (p5_y0(5),p5_y1(5),p5_y2(5),p6_y1(5),p6_y0(6));
	FA437: FA PORT MAP (p5_y0(6),p5_y1(6),p5_y2(6),p6_y1(6),p6_y0(7));
	FA438: FA PORT MAP (p5_y0(7),p5_y1(7),p5_y2(7),p6_y1(7),p6_y0(8));
	FA439: FA PORT MAP (p5_y0(8),p5_y1(8),p5_y2(8),p6_y1(8),p6_y0(9));
	FA440: FA PORT MAP (p5_y0(9),p5_y1(9),p5_y2(9),p6_y1(9),p6_y0(10));
	FA441: FA PORT MAP (p5_y0(10),p5_y1(10),p5_y2(10),p6_y1(10),p6_y0(11));
	FA442: FA PORT MAP (p5_y0(11),p5_y1(11),p5_y2(11),p6_y1(11),p6_y0(12));
	FA443: FA PORT MAP (p5_y0(12),p5_y1(12),p5_y2(12),p6_y1(12),p6_y0(13));
	FA444: FA PORT MAP (p5_y0(13),p5_y1(13),p5_y2(13),p6_y1(13),p6_y0(14));
	FA445: FA PORT MAP (p5_y0(14),p5_y1(14),p5_y2(14),p6_y1(14),p6_y0(15));
	FA446: FA PORT MAP (p5_y0(15),p5_y1(15),p5_y2(15),p6_y1(15),p6_y0(16));
	FA447: FA PORT MAP (p5_y0(16),p5_y1(16),p5_y2(16),p6_y1(16),p6_y0(17));
	FA448: FA PORT MAP (p5_y0(17),p5_y1(17),p5_y2(17),p6_y1(17),p6_y0(18));
	FA449: FA PORT MAP (p5_y0(18),p5_y1(18),p5_y2(18),p6_y1(18),p6_y0(19));
	FA450: FA PORT MAP (p5_y0(19),p5_y1(19),p5_y2(19),p6_y1(19),p6_y0(20));
	FA451: FA PORT MAP (p5_y0(20),p5_y1(20),p5_y2(20),p6_y1(20),p6_y0(21));
	FA452: FA PORT MAP (p5_y0(21),p5_y1(21),p5_y2(21),p6_y1(21),p6_y0(22));
	FA453: FA PORT MAP (p5_y0(22),p5_y1(22),p5_y2(22),p6_y1(22),p6_y0(23));
	FA454: FA PORT MAP (p5_y0(23),p5_y1(23),p5_y2(23),p6_y1(23),p6_y0(24));
	FA455: FA PORT MAP (p5_y0(24),p5_y1(24),p5_y2(24),p6_y1(24),p6_y0(25));
	FA456: FA PORT MAP (p5_y0(25),p5_y1(25),p5_y2(25),p6_y1(25),p6_y0(26));
	FA457: FA PORT MAP (p5_y0(26),p5_y1(26),p5_y2(26),p6_y1(26),p6_y0(27));
	FA458: FA PORT MAP (p5_y0(27),p5_y1(27),p5_y2(27),p6_y1(27),p6_y0(28));
	FA459: FA PORT MAP (p5_y0(28),p5_y1(28),p5_y2(28),p6_y1(28),p6_y0(29));
	FA460: FA PORT MAP (p5_y0(29),p5_y1(29),p5_y2(29),p6_y1(29),p6_y0(30));
	FA461: FA PORT MAP (p5_y0(30),p5_y1(30),p5_y2(30),p6_y1(30),p6_y0(31));
	FA462: FA PORT MAP (p5_y0(31),p5_y1(31),p5_y2(31),p6_y1(31),p6_y0(32));
	FA463: FA PORT MAP (p5_y0(32),p5_y1(32),p5_y2(32),p6_y1(32),p6_y0(33));
	FA464: FA PORT MAP (p5_y0(33),p5_y1(33),p5_y2(33),p6_y1(33),p6_y0(34));
	FA465: FA PORT MAP (p5_y0(34),p5_y1(34),p5_y2(34),p6_y1(34),p6_y0(35));
	FA466: FA PORT MAP (p5_y0(35),p5_y1(35),p5_y2(35),p6_y1(35),p6_y0(36));
	FA467: FA PORT MAP (p5_y0(36),p5_y1(36),p5_y2(36),p6_y1(36),p6_y0(37));
	FA468: FA PORT MAP (p5_y0(37),p5_y1(37),p5_y2(37),p6_y1(37),p6_y0(38));
	FA469: FA PORT MAP (p5_y0(38),p5_y1(38),p5_y2(38),p6_y1(38),p6_y0(39));
	FA470: FA PORT MAP (p5_y0(39),p5_y1(39),p5_y2(39),p6_y1(39),p6_y0(40));
	FA471: FA PORT MAP (p5_y0(40),p5_y1(40),p5_y2(40),p6_y1(40),p6_y0(41));
	FA472: FA PORT MAP (p5_y0(41),p5_y1(41),p5_y2(41),p6_y1(41),p6_y0(42));
	FA473: FA PORT MAP (p5_y0(42),p5_y1(42),p5_y2(42),p6_y1(42),p6_y0(43));
	FA474: FA PORT MAP (p5_y0(43),p5_y1(43),p5_y2(43),p6_y1(43),p6_y0(44));
	FA475: FA PORT MAP (p5_y0(44),p5_y1(44),p5_y2(44),p6_y1(44),p6_y0(45));
	FA476: FA PORT MAP (p5_y0(45),p5_y1(45),p5_y2(45),p6_y1(45),p6_y0(46));
	FA477: FA PORT MAP (p5_y0(46),p5_y1(46),p5_y2(46),p6_y1(46),p6_y0(47));
	FA478: FA PORT MAP (p5_y0(47),p5_y1(47),p5_y2(47),p6_y1(47),p6_y0(48));
	FA479: FA PORT MAP (p5_y0(48),p5_y1(48),p5_y2(48),p6_y1(48),p6_y0(49));
	FA480: FA PORT MAP (p5_y0(49),p5_y1(49),p5_y2(49),p6_y1(49),p6_y0(50));
	FA481: FA PORT MAP (p5_y0(50),p5_y1(50),p5_y2(50),p6_y1(50),p6_y0(51));
	FA482: FA PORT MAP (p5_y0(51),p5_y1(51),p5_y2(51),p6_y1(51),p6_y0(52));
	FA483: FA PORT MAP (p5_y0(52),p5_y1(52),p5_y2(52),p6_y1(52),p6_y0(53));
	FA484: FA PORT MAP (p5_y0(53),p5_y1(53),p5_y2(53),p6_y1(53),p6_y0(54));
	FA485: FA PORT MAP (p5_y0(54),p5_y1(54),p5_y2(54),p6_y1(54),p6_y0(55));
	FA486: FA PORT MAP (p5_y0(55),p5_y1(55),p5_y2(55),p6_y1(55),p6_y0(56));
	FA487: FA PORT MAP (p5_y0(56),p5_y1(56),p5_y2(56),p6_y1(56),p6_y0(57));
	FA488: FA PORT MAP (p5_y0(57),p5_y1(57),p5_y2(57),p6_y1(57),p6_y0(58));
	FA489: FA PORT MAP (p5_y0(58),p5_y1(58),p5_y2(58),p6_y1(58),p6_y0(59));
	FA490: FA PORT MAP (p5_y0(59),p5_y1(59),p5_y2(59),p6_y1(59),p6_y0(60));
	FA491: FA PORT MAP (p5_y0(60),p5_y1(60),p5_y2(60),p6_y1(60),p6_y0(61));
	FA492: FA PORT MAP (p5_y0(61),p5_y1(61),p5_y2(61),p6_y1(61),p6_y0(62));
	FA493: FA PORT MAP (p5_y0(62),p5_y1(62),p5_y2(62),p6_y1(62),p6_y0(63));
	FA494: FA PORT MAP (p5_y0(63),p5_y1(63),p5_y2(63),p6_y1(63),overflow_bit);
	
	product <= std_logic_vector(unsigned(p6_y1)+unsigned(p6_y0));
	
end beh;

