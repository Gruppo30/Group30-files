LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.ALL;

entity regFile is
	generic (  k : positive := 5;
               N : integer := 64);
	port(	clock,rst : in std_logic;
			rs1	 	  : in  unsigned ((k-1) downto 0);
			rs2		  : in  unsigned ((k-1) downto 0);
			rd 		  : in  unsigned ((k-1) downto 0);
			data_in   : in  std_logic_vector ((N-1) downto 0);
			wr_en	  : in  std_logic;
			data1_out : out std_logic_vector ((N-1) downto 0);
			data2_out : out std_logic_vector ((N-1) downto 0)
		);
end regFile;

architecture beh of regFile is

	signal data_in_tmp : std_logic_vector ((N-1) downto 0);

	type regF is array(0 to (2**k)-1) of std_logic_vector ((N-1) downto 0);
	signal regArray : regF;
	

begin 
	
	
	process(rs1, rs2, clock, rst, wr_en, rd, data_in, regArray)
	begin
		if (rst = '0') then
				regArray <= (	"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000",
								"0000000000000000000000000000000000000000000000000000000000000000");
			data1_out <= (others => '0');
			data2_out <= (others => '0');		
			
		else 
		if((rs1=rd) and (wr_en='1'))then data1_out<=data_in;
		else data1_out <= regArray(to_integer(rs1)); end if;
	
		if((rs2=rd) and (wr_en='1'))then data2_out<=data_in;
		else data2_out <= regArray(to_integer(rs2)); end if;
		
		if(clock'event and clock='1' and wr_en = '1') then
			regArray(to_integer(rd)) <= data_in;
		end if;
		end if;
		
	end process;
end beh;
